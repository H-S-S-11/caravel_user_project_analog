magic
tech sky130A
magscale 1 2
timestamp 1635946216
<< error_p >>
rect 3831 2230 3871 2266
rect 3835 2148 3871 2230
rect 3831 2112 3871 2148
rect 3861 1845 3895 1847
rect 3861 1829 3895 1831
rect 3861 1791 3895 1793
rect 3861 1777 3895 1779
rect 3861 1757 3895 1759
rect 3861 1719 3895 1721
rect 3861 1709 3895 1711
rect 3861 1685 3895 1687
rect 3861 1647 3895 1649
rect 3861 1641 3895 1643
rect 3861 1613 3895 1615
rect 3861 1573 3895 1577
rect 3861 1541 3895 1543
rect 3861 1503 3895 1507
rect 3861 1469 3895 1471
rect 3861 1437 3895 1439
rect 3861 1431 3895 1433
rect 3861 1397 3895 1399
rect 3861 1369 3895 1371
rect 3861 1359 3895 1361
rect 3861 1325 3895 1327
rect 3861 1301 3895 1303
rect 3861 1287 3895 1289
rect 3861 1253 3895 1255
rect 3861 1233 3895 1235
rect 3861 1215 3895 1217
rect 3861 1181 3895 1183
rect 3861 1165 3895 1167
rect 3861 1143 3895 1145
rect 3861 1109 3895 1111
rect 3861 1097 3895 1099
rect 3861 1071 3895 1073
rect 3861 1037 3895 1039
rect 3861 1029 3895 1031
rect 3861 999 3895 1001
rect 3861 965 3895 967
rect 3861 961 3895 963
rect 3861 927 3895 929
rect 3861 893 3895 895
rect 3861 855 3895 857
rect 3861 825 3895 827
rect 3861 821 3895 823
rect 3861 783 3895 785
rect 3861 757 3895 759
rect 3861 749 3895 751
rect 3861 711 3895 713
rect 3861 689 3895 691
rect 3861 677 3895 679
rect 3861 639 3895 641
rect 3861 621 3895 623
rect 3861 605 3895 607
rect 3861 567 3895 569
rect 3861 553 3895 555
rect 3861 533 3895 535
rect 3861 495 3895 497
rect 3861 485 3895 487
rect 3861 461 3895 463
rect 3861 423 3895 425
rect 3861 417 3895 419
rect 3861 389 3895 391
rect 3861 349 3895 353
rect 3861 317 3895 319
rect 3861 279 3895 283
rect 3861 245 3895 247
rect 3861 213 3895 215
rect 3861 207 3895 209
rect 3861 173 3895 175
rect 3861 145 3895 147
rect 3861 135 3895 137
rect 3861 101 3895 103
rect 3861 77 3895 79
rect 3861 63 3895 65
rect 3861 29 3895 31
rect 3861 9 3895 11
rect 3861 -9 3895 -7
use m10_nfet_w10_l1  m10_nfet_w10_l1_0
array 0 1 8000 0 0 0
timestamp 1635946216
transform 1 0 -197 0 1 18
box -2712 -817 4234 2603
<< end >>
