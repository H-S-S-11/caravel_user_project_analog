magic
tech sky130A
magscale 1 2
timestamp 1632403905
<< pwell >>
rect -214 -1146 214 1146
<< nmos >>
rect -18 736 18 936
rect -18 318 18 518
rect -18 -100 18 100
rect -18 -518 18 -318
rect -18 -936 18 -736
<< ndiff >>
rect -76 924 -18 936
rect -76 748 -64 924
rect -30 748 -18 924
rect -76 736 -18 748
rect 18 924 76 936
rect 18 748 30 924
rect 64 748 76 924
rect 18 736 76 748
rect -76 506 -18 518
rect -76 330 -64 506
rect -30 330 -18 506
rect -76 318 -18 330
rect 18 506 76 518
rect 18 330 30 506
rect 64 330 76 506
rect 18 318 76 330
rect -76 88 -18 100
rect -76 -88 -64 88
rect -30 -88 -18 88
rect -76 -100 -18 -88
rect 18 88 76 100
rect 18 -88 30 88
rect 64 -88 76 88
rect 18 -100 76 -88
rect -76 -330 -18 -318
rect -76 -506 -64 -330
rect -30 -506 -18 -330
rect -76 -518 -18 -506
rect 18 -330 76 -318
rect 18 -506 30 -330
rect 64 -506 76 -330
rect 18 -518 76 -506
rect -76 -748 -18 -736
rect -76 -924 -64 -748
rect -30 -924 -18 -748
rect -76 -936 -18 -924
rect 18 -748 76 -736
rect 18 -924 30 -748
rect 64 -924 76 -748
rect 18 -936 76 -924
<< ndiffc >>
rect -64 748 -30 924
rect 30 748 64 924
rect -64 330 -30 506
rect 30 330 64 506
rect -64 -88 -30 88
rect 30 -88 64 88
rect -64 -506 -30 -330
rect 30 -506 64 -330
rect -64 -924 -30 -748
rect 30 -924 64 -748
<< psubdiff >>
rect -178 1076 -82 1110
rect 82 1076 178 1110
rect -178 1014 -144 1076
rect 144 1014 178 1076
rect -178 -583 -144 537
rect -178 -1076 -144 -1014
rect 144 -1076 178 -1014
rect -178 -1110 -82 -1076
rect 82 -1110 178 -1076
<< psubdiffcont >>
rect -82 1076 82 1110
rect -178 537 -144 1014
rect -178 -1014 -144 -583
rect 144 -1014 178 1014
rect -82 -1110 82 -1076
<< poly >>
rect -33 1008 33 1024
rect -33 974 -17 1008
rect 17 974 33 1008
rect -33 958 33 974
rect -18 936 18 958
rect -18 714 18 736
rect -33 698 33 714
rect -33 664 -17 698
rect 17 664 33 698
rect -33 648 33 664
rect -33 590 33 606
rect -33 556 -17 590
rect 17 556 33 590
rect -33 540 33 556
rect -18 518 18 540
rect -18 296 18 318
rect -33 280 33 296
rect -33 246 -17 280
rect 17 246 33 280
rect -33 230 33 246
rect -33 172 33 188
rect -33 138 -17 172
rect 17 138 33 172
rect -33 122 33 138
rect -18 100 18 122
rect -18 -122 18 -100
rect -33 -138 33 -122
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -33 -188 33 -172
rect -33 -246 33 -230
rect -33 -280 -17 -246
rect 17 -280 33 -246
rect -33 -296 33 -280
rect -18 -318 18 -296
rect -18 -540 18 -518
rect -33 -556 33 -540
rect -33 -590 -17 -556
rect 17 -590 33 -556
rect -33 -606 33 -590
rect -33 -664 33 -648
rect -33 -698 -17 -664
rect 17 -698 33 -664
rect -33 -714 33 -698
rect -18 -736 18 -714
rect -18 -958 18 -936
rect -33 -974 33 -958
rect -33 -1008 -17 -974
rect 17 -1008 33 -974
rect -33 -1024 33 -1008
<< polycont >>
rect -17 974 17 1008
rect -17 664 17 698
rect -17 556 17 590
rect -17 246 17 280
rect -17 138 17 172
rect -17 -172 17 -138
rect -17 -280 17 -246
rect -17 -590 17 -556
rect -17 -698 17 -664
rect -17 -1008 17 -974
<< locali >>
rect -178 1076 -82 1110
rect 82 1076 178 1110
rect -178 1014 -144 1076
rect -201 537 -178 567
rect 144 1014 178 1076
rect -33 974 -17 1008
rect 17 974 33 1008
rect -64 924 -30 940
rect -64 732 -30 748
rect 30 924 64 940
rect 30 732 64 748
rect -33 664 -17 698
rect 17 664 33 698
rect -144 537 -121 567
rect -33 556 -17 590
rect 17 556 33 590
rect -201 517 -121 537
rect -64 506 -30 522
rect -64 314 -30 330
rect 30 506 64 522
rect 30 314 64 330
rect -33 246 -17 280
rect 17 246 33 280
rect -33 138 -17 172
rect 17 138 33 172
rect -64 88 -30 104
rect -64 -104 -30 -88
rect 30 88 64 104
rect 30 -104 64 -88
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -33 -280 -17 -246
rect 17 -280 33 -246
rect -64 -330 -30 -314
rect -64 -522 -30 -506
rect 30 -330 64 -314
rect 30 -522 64 -506
rect -201 -583 -121 -563
rect -201 -603 -178 -583
rect -144 -603 -121 -583
rect -33 -590 -17 -556
rect 17 -590 33 -556
rect -33 -698 -17 -664
rect 17 -698 33 -664
rect -64 -748 -30 -732
rect -64 -940 -30 -924
rect 30 -748 64 -732
rect 30 -940 64 -924
rect -33 -1008 -17 -974
rect 17 -1008 33 -974
rect -178 -1076 -144 -1014
rect 144 -1076 178 -1014
rect -178 -1110 -82 -1076
rect 82 -1110 178 -1076
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -161 -1093 161 1093
string parameters w 1 l 0.18 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
