magic
tech sky130A
timestamp 1634766604
<< nwell >>
rect 1400 -2600 1900 -2100
<< nnmos >>
rect 980 -2240 1050 -2190
rect 980 -2370 1050 -2320
rect 980 -2480 1050 -2430
<< mvpmos >>
rect 1500 -2240 1600 -2190
rect 1500 -2370 1600 -2320
rect 1500 -2480 1600 -2430
<< mvndiff >>
rect 980 -2160 1050 -2150
rect 980 -2180 990 -2160
rect 1040 -2180 1050 -2160
rect 980 -2190 1050 -2180
rect 980 -2250 1050 -2240
rect 980 -2310 990 -2250
rect 1040 -2310 1050 -2250
rect 980 -2320 1050 -2310
rect 980 -2430 1050 -2370
rect 980 -2490 1050 -2480
rect 980 -2510 990 -2490
rect 1040 -2510 1050 -2490
rect 980 -2520 1050 -2510
<< mvpdiff >>
rect 1500 -2160 1600 -2150
rect 1500 -2180 1510 -2160
rect 1590 -2180 1600 -2160
rect 1500 -2190 1600 -2180
rect 1500 -2250 1600 -2240
rect 1500 -2310 1510 -2250
rect 1590 -2310 1600 -2250
rect 1500 -2320 1600 -2310
rect 1500 -2380 1600 -2370
rect 1500 -2410 1510 -2380
rect 1590 -2410 1600 -2380
rect 1500 -2430 1600 -2410
rect 1500 -2490 1600 -2480
rect 1500 -2510 1510 -2490
rect 1590 -2510 1600 -2490
rect 1500 -2520 1600 -2510
<< mvndiffc >>
rect 990 -2180 1040 -2160
rect 990 -2310 1040 -2250
rect 990 -2510 1040 -2490
<< mvpdiffc >>
rect 1510 -2180 1590 -2160
rect 1510 -2310 1590 -2250
rect 1510 -2410 1590 -2380
rect 1510 -2510 1590 -2490
<< poly >>
rect 1220 -2190 1340 -2180
rect 960 -2240 980 -2190
rect 1050 -2240 1230 -2190
rect 1330 -2240 1500 -2190
rect 1600 -2240 1620 -2190
rect 1220 -2250 1340 -2240
rect 960 -2370 980 -2320
rect 1050 -2370 1500 -2320
rect 1600 -2370 1620 -2320
rect 960 -2480 980 -2430
rect 1050 -2480 1500 -2430
rect 1600 -2480 1620 -2430
<< polycont >>
rect 1230 -2240 1330 -2190
<< locali >>
rect 800 1850 1050 1900
rect 1500 1850 1750 1900
rect 800 -1950 1050 -1900
rect 980 -2100 1050 -1950
rect 1500 -1950 1750 -1900
rect 1500 -1970 1550 -1950
rect 980 -2160 1050 -2150
rect 980 -2180 990 -2160
rect 1040 -2180 1050 -2160
rect 1400 -2020 1550 -1970
rect 1220 -2190 1340 -2180
rect 1400 -2190 1450 -2020
rect 1500 -2160 1600 -2150
rect 1500 -2180 1510 -2160
rect 1590 -2180 1600 -2160
rect 1100 -2240 1230 -2190
rect 1330 -2240 1450 -2190
rect 790 -2310 990 -2250
rect 1040 -2310 1050 -2250
rect 1100 -2490 1150 -2240
rect 1220 -2250 1340 -2240
rect 1400 -2380 1450 -2240
rect 1500 -2310 1510 -2250
rect 1590 -2310 1790 -2250
rect 1400 -2410 1510 -2380
rect 1590 -2410 1600 -2380
rect 980 -2510 990 -2490
rect 1040 -2510 1150 -2490
rect 980 -2520 1150 -2510
rect 1500 -2510 1510 -2490
rect 1590 -2510 1790 -2490
rect 1500 -2520 1790 -2510
<< viali >>
rect 980 -2150 1050 -2100
rect 1500 -2150 1600 -2100
<< metal1 >>
rect 2750 1150 2800 1550
rect -50 350 0 750
rect 2750 -750 2800 -350
rect -50 -1550 0 -1150
rect 970 -2100 1610 -2090
rect 970 -2150 980 -2100
rect 1050 -2150 1500 -2100
rect 1600 -2150 1610 -2100
rect 970 -2160 1610 -2150
<< metal2 >>
rect 100 1850 600 1900
rect 2150 1850 2650 1900
rect 100 -50 600 0
rect 2150 -50 2650 0
rect 100 -1950 600 -1900
rect 2150 -1950 2650 -1900
use analog_switch  analog_switch_1
timestamp 1634419951
transform 1 0 500 0 1 -1150
box -500 -750 2250 1100
use analog_switch  analog_switch_0
timestamp 1634419951
transform 1 0 500 0 1 750
box -500 -750 2250 1100
<< labels >>
rlabel locali 990 -2040 1040 -1990 1 EN0
rlabel locali 1450 -2010 1490 -1980 1 ENB0
<< end >>
