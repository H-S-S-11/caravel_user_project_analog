magic
tech sky130A
magscale 1 2
timestamp 1635946216
<< pwell >>
rect -103 -67 103 67
<< locali >>
rect -69 -33 69 33
<< end >>
