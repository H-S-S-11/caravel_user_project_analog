magic
tech sky130A
magscale 1 2
timestamp 1632245862
<< nwell >>
rect 60 1210 150 1540
rect 0 1170 150 1210
rect 0 1060 150 1100
rect 60 730 150 1060
<< pwell >>
rect 880 1260 950 1440
rect 620 1160 850 1210
rect 620 1070 850 1120
rect 890 840 950 1020
rect 660 330 910 460
<< locali >>
rect -80 2440 180 2460
rect -80 2340 -60 2440
rect 160 2340 180 2440
rect -80 2280 180 2340
rect 640 2200 920 2220
rect -160 1780 270 2170
rect 640 2100 660 2200
rect 900 2100 920 2200
rect 640 2040 920 2100
rect 1300 2000 1760 2020
rect 660 1860 910 1950
rect 1300 1900 1320 2000
rect 1740 1900 1760 2000
rect 550 1820 1010 1860
rect 1300 1840 1760 1900
rect 550 1680 700 1820
rect 860 1680 1010 1820
rect 1460 1750 1610 1840
rect 1330 1660 1730 1750
rect -160 1260 -20 1540
rect 60 1440 150 1540
rect 1220 1480 1850 1660
rect 60 1210 150 1350
rect 1330 1390 1730 1480
rect 0 1170 150 1210
rect 660 1170 850 1210
rect 620 1160 850 1170
rect 620 1110 850 1120
rect 0 1060 150 1100
rect 660 1070 850 1110
rect 1220 1080 1360 1240
rect 1490 1180 1570 1190
rect 1490 1120 1500 1180
rect 1560 1120 1570 1180
rect 1490 1110 1570 1120
rect 1210 1070 1360 1080
rect 1700 1080 1840 1240
rect 1700 1070 1850 1080
rect 1210 1060 1350 1070
rect 1710 1060 1850 1070
rect -160 730 -20 1010
rect 60 930 150 1060
rect 60 730 150 840
rect 1330 820 1730 910
rect 1220 640 1840 820
rect -160 100 270 490
rect 550 460 700 600
rect 860 460 1010 600
rect 1330 550 1730 640
rect 550 420 1010 460
rect 1460 440 1610 550
rect 660 330 910 420
<< viali >>
rect -60 2340 160 2440
rect 660 2100 900 2200
rect 1320 1900 1740 2000
rect 60 1350 150 1440
rect 630 1350 690 1440
rect 860 1260 950 1440
rect 1400 1290 1490 1330
rect 1580 1290 1670 1330
rect 620 1170 660 1210
rect 620 1070 660 1110
rect 1500 1120 1560 1180
rect 60 840 150 930
rect 630 840 690 930
rect 860 840 950 1020
<< metal1 >>
rect -80 2440 180 2460
rect -80 2340 -60 2440
rect 160 2340 180 2440
rect -80 2320 180 2340
rect 640 2200 1760 2460
rect 640 2100 660 2200
rect 900 2100 1760 2200
rect 640 2080 1760 2100
rect 1300 2000 1760 2080
rect 1300 1900 1320 2000
rect 1740 1900 1760 2000
rect 1300 1880 1760 1900
rect 40 1440 710 1460
rect 40 1350 60 1440
rect 150 1350 630 1440
rect 690 1350 710 1440
rect 40 1330 710 1350
rect 840 1440 970 1460
rect 840 1260 860 1440
rect 950 1260 970 1440
rect 1380 1330 1690 1350
rect 1380 1290 1400 1330
rect 1490 1290 1580 1330
rect 1670 1290 1690 1330
rect 1380 1270 1690 1290
rect 600 1210 680 1230
rect 600 1170 620 1210
rect 660 1170 680 1210
rect 600 1160 680 1170
rect 840 1200 970 1260
rect 840 1180 1580 1200
rect 840 1120 1500 1180
rect 1560 1120 1580 1180
rect 600 1110 680 1120
rect 600 1070 620 1110
rect 660 1070 680 1110
rect 600 1050 680 1070
rect 840 1100 1580 1120
rect 840 1020 970 1100
rect 40 930 710 950
rect 40 840 60 930
rect 150 840 630 930
rect 690 840 710 930
rect 40 820 710 840
rect 840 840 860 1020
rect 950 840 970 1020
rect 840 820 970 840
use sky130_fd_pr__nfet_03v3_nvt_DWHJCV  sky130_fd_pr__nfet_03v3_nvt_DWHJCV_0
timestamp 1632244313
transform 1 0 1532 0 1 1151
box -377 -776 377 776
use sky130_fd_pr__nfet_03v3_nvt_ZJHJCF  sky130_fd_pr__nfet_03v3_nvt_ZJHJCF_0
timestamp 1632244518
transform 1 0 783 0 1 1140
box -288 -985 288 985
use sky130_fd_pr__pfet_g5v0d10v5_CABTE7  sky130_fd_pr__pfet_g5v0d10v5_CABTE7_0
timestamp 1632243750
transform 1 0 53 0 1 1136
box -308 -1251 308 1251
<< labels >>
rlabel metal1 640 2380 1760 2460 1 VGND
rlabel metal1 -80 2420 180 2460 1 VPWR
rlabel metal1 1480 1100 1580 1200 1 VI
rlabel metal1 1380 1270 1690 1350 1 BIASN
rlabel metal1 390 1330 460 1460 1 VPAMP
rlabel metal1 390 820 460 950 1 VNAMP
rlabel metal1 600 1160 680 1230 1 VP
rlabel metal1 600 1050 680 1120 1 VN
<< end >>
