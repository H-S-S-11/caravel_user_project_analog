magic
tech sky130A
magscale 1 4
timestamp 1632405528
<< nwell >>
rect -880 5200 1240 6200
rect -40 2280 1240 5200
<< pwell >>
rect -1840 5040 -960 6560
rect -1840 4000 -320 5040
rect -1840 1960 -960 4000
<< nmos >>
rect -640 4560 -580 4960
<< pmos >>
rect -640 5280 -580 6080
<< ndiff >>
rect -800 4920 -640 4960
rect -800 4600 -760 4920
rect -680 4600 -640 4920
rect -800 4560 -640 4600
rect -580 4920 -400 4960
rect -580 4600 -520 4920
rect -440 4600 -400 4920
rect -580 4560 -400 4600
<< pdiff >>
rect -800 6040 -640 6080
rect -800 5320 -760 6040
rect -680 5320 -640 6040
rect -800 5280 -640 5320
rect -580 6040 -400 6080
rect -580 5320 -520 6040
rect -440 5320 -400 6040
rect -580 5280 -400 5320
<< ndiffc >>
rect -760 4600 -680 4920
rect -520 4600 -440 4920
<< pdiffc >>
rect -760 5320 -680 6040
rect -520 5320 -440 6040
<< psubdiff >>
rect -640 4360 -360 4440
rect -640 4240 -560 4360
rect -440 4240 -360 4360
rect -640 4160 -360 4240
<< psubdiffcont >>
rect -560 4240 -440 4360
<< poly >>
rect -640 6080 -580 6140
rect -640 5160 -580 5280
rect -320 5160 -120 5200
rect -640 5040 -280 5160
rect -160 5040 -120 5160
rect -640 4960 -580 5040
rect -320 5000 -120 5040
rect -640 4490 -580 4560
<< polycont >>
rect -280 5040 -160 5160
<< locali >>
rect -1720 5640 -1080 6440
rect -800 6360 -520 6480
rect -800 6040 -680 6360
rect -800 5320 -760 6040
rect -1760 5040 -1480 5200
rect -1760 4360 -1640 5040
rect -800 4920 -680 5320
rect -520 6040 280 6080
rect 960 6040 1120 6080
rect -440 5320 1120 6040
rect -520 5280 1120 5320
rect 120 5240 1120 5280
rect -320 5160 -120 5200
rect -320 5040 -280 5160
rect -160 5040 -120 5160
rect -320 5000 -120 5040
rect 480 4980 1140 5060
rect -800 4600 -760 4920
rect -800 4560 -680 4600
rect -520 4920 -400 4960
rect -440 4600 -400 4920
rect -520 4440 -400 4600
rect -640 4400 -360 4440
rect -1760 4200 -1480 4360
rect -1760 3520 -1640 4200
rect -1320 4160 -1080 4360
rect -640 4200 -600 4400
rect -400 4200 -360 4400
rect 280 4340 380 4960
rect 480 4460 560 4980
rect 660 4340 760 4900
rect 860 4460 940 4980
rect 280 4260 760 4340
rect -640 4160 -360 4200
rect 480 4100 1100 4180
rect -1400 3900 -1320 3980
rect -1480 3780 -1380 3800
rect -1480 3720 -1340 3780
rect 240 3520 380 4020
rect 480 3600 560 4100
rect 660 3520 760 4020
rect 860 3580 940 4100
rect -1760 3360 -1520 3520
rect 240 3480 760 3520
rect 360 3420 760 3480
rect -1720 2080 -1080 2880
rect 120 2400 1120 3240
<< viali >>
rect -1560 6440 -1240 6720
rect -520 6360 -400 6480
rect -1080 5360 -880 5560
rect -1320 5000 -1240 5200
rect 280 6040 960 6440
rect -280 5040 -160 5160
rect 240 4960 400 5160
rect -1440 4740 -1360 4820
rect -1080 4640 -880 4840
rect -600 4360 -400 4400
rect -600 4240 -560 4360
rect -560 4240 -440 4360
rect -440 4240 -400 4360
rect -600 4200 -400 4240
rect -1320 3900 -1240 3980
rect -1560 3720 -1480 3800
rect -1320 3320 -1240 3520
rect 240 3360 360 3480
<< metal1 >>
rect -1600 6720 -840 6800
rect -1600 6440 -1560 6720
rect -1240 6440 -840 6720
rect -1600 6400 -840 6440
rect -1120 5560 -840 6400
rect -560 6480 -360 6800
rect -560 6360 -520 6480
rect -400 6360 -360 6480
rect -560 6320 -360 6360
rect 200 6440 1040 6800
rect 200 6040 280 6440
rect 960 6040 1040 6440
rect 200 5960 1040 6040
rect -1120 5360 -1080 5560
rect -880 5360 -840 5560
rect -1120 5320 -840 5360
rect -1360 5200 -1200 5240
rect -1360 5000 -1320 5200
rect -1240 5160 -1200 5200
rect -320 5160 -120 5200
rect 200 5160 440 5200
rect -1240 5040 -280 5160
rect -160 5040 240 5160
rect -1240 5000 -1200 5040
rect -320 5000 -120 5040
rect -1360 4960 -1200 5000
rect 200 4960 240 5040
rect 400 4960 440 5160
rect 200 4920 440 4960
rect -1120 4840 -840 4880
rect -1880 4820 -1320 4840
rect -1880 4740 -1440 4820
rect -1360 4740 -1320 4820
rect -1880 4720 -1320 4740
rect -1120 4640 -1080 4840
rect -880 4640 -840 4840
rect -1120 4440 -840 4640
rect -1120 4400 -360 4440
rect -1120 4200 -600 4400
rect -400 4200 -360 4400
rect -1120 4160 -360 4200
rect -1360 3980 -1200 4020
rect -1360 3900 -1320 3980
rect -1240 3900 -1200 3980
rect -1360 3860 -1200 3900
rect -1880 3800 -1440 3840
rect -1880 3720 -1560 3800
rect -1480 3720 -1440 3800
rect -1600 3680 -1440 3720
rect -1320 3560 -1240 3860
rect -1360 3520 -1200 3560
rect -1360 3320 -1320 3520
rect -1240 3480 -1200 3520
rect 200 3480 400 3520
rect -1240 3360 240 3480
rect 360 3360 400 3480
rect -1240 3320 -1200 3360
rect 200 3320 400 3360
rect -1360 3280 -1200 3320
use sky130_fd_pr__nfet_01v8_T49HPK  sky130_fd_pr__nfet_01v8_T49HPK_0
timestamp 1632403905
transform 1 0 -1398 0 1 4266
box -428 -2292 428 2292
use sky130_fd_pr__pfet_01v8_XAY5ZQ  sky130_fd_pr__pfet_01v8_XAY5ZQ_0
timestamp 1632400215
transform 1 0 613 0 1 4240
box -619 -1946 619 1946
<< labels >>
rlabel metal1 200 6760 1040 6800 1 VPWR
rlabel locali -1640 5080 -1560 5160 1 ISINK
rlabel metal1 -1880 3720 -1840 3840 1 VON
rlabel metal1 -1880 4720 -1840 4840 1 VOP
rlabel metal1 -920 5040 -840 5160 1 VOPAMP
rlabel metal1 -840 3360 -720 3480 1 VONAMP
rlabel metal1 -1600 6760 -840 6800 1 VGND
rlabel metal1 -560 6760 -360 6800 1 VOUT
<< end >>
