magic
tech sky130A
timestamp 1633173629
<< pwell >>
rect -80 -50 80 210
<< nnmos >>
rect -30 90 20 190
rect -25 -21 25 21
<< mvndiff >>
rect -70 180 -30 190
rect -70 100 -60 180
rect -40 100 -30 180
rect -70 90 -30 100
rect 20 180 60 190
rect 20 100 30 180
rect 50 100 60 180
rect 20 90 60 100
rect -55 15 -25 21
rect -55 -15 -49 15
rect -31 -15 -25 15
rect -55 -21 -25 -15
rect 25 15 55 21
rect 25 -15 31 15
rect 49 -15 55 15
rect 25 -21 55 -15
<< mvndiffc >>
rect -60 100 -40 180
rect 30 100 50 180
rect -49 -15 -31 15
rect 31 -15 49 15
<< poly >>
rect -30 190 20 210
rect -30 70 20 90
rect -25 21 25 34
rect -25 -34 25 -21
<< locali >>
rect -70 180 -40 190
rect -70 100 -60 180
rect -70 90 -40 100
rect 30 180 60 190
rect 50 100 60 180
rect 30 90 60 100
rect -50 15 -30 30
rect -50 -15 -49 15
rect -31 -15 -30 15
rect -50 -30 -30 -15
rect 30 15 50 30
rect 30 -15 31 15
rect 49 -15 50 15
rect 30 -30 50 -15
<< end >>
