magic
tech sky130A
magscale 1 2
timestamp 1632242116
<< nwell >>
rect -308 -1251 308 1251
<< mvpmos >>
rect -50 654 50 954
rect -50 118 50 418
rect -50 -418 50 -118
rect -50 -954 50 -654
<< mvpdiff >>
rect -108 942 -50 954
rect -108 666 -96 942
rect -62 666 -50 942
rect -108 654 -50 666
rect 50 942 108 954
rect 50 666 62 942
rect 96 666 108 942
rect 50 654 108 666
rect -108 406 -50 418
rect -108 130 -96 406
rect -62 130 -50 406
rect -108 118 -50 130
rect 50 406 108 418
rect 50 130 62 406
rect 96 130 108 406
rect 50 118 108 130
rect -108 -130 -50 -118
rect -108 -406 -96 -130
rect -62 -406 -50 -130
rect -108 -418 -50 -406
rect 50 -130 108 -118
rect 50 -406 62 -130
rect 96 -406 108 -130
rect 50 -418 108 -406
rect -108 -666 -50 -654
rect -108 -942 -96 -666
rect -62 -942 -50 -666
rect -108 -954 -50 -942
rect 50 -666 108 -654
rect 50 -942 62 -666
rect 96 -942 108 -666
rect 50 -954 108 -942
<< mvpdiffc >>
rect -96 666 -62 942
rect 62 666 96 942
rect -96 130 -62 406
rect 62 130 96 406
rect -96 -406 -62 -130
rect 62 -406 96 -130
rect -96 -942 -62 -666
rect 62 -942 96 -666
<< mvnsubdiff >>
rect -242 1173 242 1185
rect -242 1139 -134 1173
rect 134 1139 242 1173
rect -242 1127 242 1139
rect -242 1077 -184 1127
rect -242 -1077 -230 1077
rect -196 -1077 -184 1077
rect 184 1077 242 1127
rect -242 -1127 -184 -1077
rect 184 -1077 196 1077
rect 230 -1077 242 1077
rect 184 -1127 242 -1077
rect -242 -1139 242 -1127
rect -242 -1173 -134 -1139
rect 134 -1173 242 -1139
rect -242 -1185 242 -1173
<< mvnsubdiffcont >>
rect -134 1139 134 1173
rect -230 -1077 -196 1077
rect 196 -1077 230 1077
rect -134 -1173 134 -1139
<< poly >>
rect -50 1035 50 1051
rect -50 1001 -34 1035
rect 34 1001 50 1035
rect -50 954 50 1001
rect -50 607 50 654
rect -50 573 -34 607
rect 34 573 50 607
rect -50 557 50 573
rect -50 499 50 515
rect -50 465 -34 499
rect 34 465 50 499
rect -50 418 50 465
rect -50 71 50 118
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -118 50 -71
rect -50 -465 50 -418
rect -50 -499 -34 -465
rect 34 -499 50 -465
rect -50 -515 50 -499
rect -50 -573 50 -557
rect -50 -607 -34 -573
rect 34 -607 50 -573
rect -50 -654 50 -607
rect -50 -1001 50 -954
rect -50 -1035 -34 -1001
rect 34 -1035 50 -1001
rect -50 -1051 50 -1035
<< polycont >>
rect -34 1001 34 1035
rect -34 573 34 607
rect -34 465 34 499
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -499 34 -465
rect -34 -607 34 -573
rect -34 -1035 34 -1001
<< locali >>
rect -230 1139 -134 1173
rect 134 1139 230 1173
rect -230 1077 -196 1139
rect 196 1077 230 1139
rect -50 1001 -34 1035
rect 34 1001 50 1035
rect -96 942 -62 958
rect -96 650 -62 666
rect 62 942 96 958
rect 62 650 96 666
rect -50 573 -34 607
rect 34 573 50 607
rect -50 465 -34 499
rect 34 465 50 499
rect -96 406 -62 422
rect -96 114 -62 130
rect 62 406 96 422
rect 62 114 96 130
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -130 -62 -114
rect -96 -422 -62 -406
rect 62 -130 96 -114
rect 62 -422 96 -406
rect -50 -499 -34 -465
rect 34 -499 50 -465
rect -50 -607 -34 -573
rect 34 -607 50 -573
rect -96 -666 -62 -650
rect -96 -958 -62 -942
rect 62 -666 96 -650
rect 62 -958 96 -942
rect -50 -1035 -34 -1001
rect 34 -1035 50 -1001
rect -230 -1139 -196 -1077
rect 196 -1139 230 -1077
rect -230 -1173 -134 -1139
rect 134 -1173 230 -1139
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string FIXED_BBOX -213 -1156 213 1156
string parameters w 1.5 l 0.5 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
