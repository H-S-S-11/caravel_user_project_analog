**.subckt chargepump_tb
x1 VIN vout VCLK chargepump
V1 VIN GND 3
V2 VCLK GND PULSE(0 3 100n 1n 1n 100n 200n)
**** begin user architecture code


.lib ~/open_sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt


.control
tran 10n 100u
plot V(VIN) V(vout) v(VCLK)
.endc

**** end user architecture code
**.ends

* expanding   symbol:  chargepump.sym # of pins=3
* sym_path: /home/hss11/winhome/skywater-shuttle/caravel_user_project_analog/xschem/chargepump.sym
* sch_path: /home/hss11/winhome/skywater-shuttle/caravel_user_project_analog/xschem/chargepump.sch
.subckt chargepump  VIN VOUT CLKIN
*.ipin VIN
*.ipin CLKIN
*.opin VOUT
XM2 VOUT net1 net1 net1 sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 VOUT net1 net1 net1 sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 net1 VIN VIN VIN sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 net1 VIN VIN VIN sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XC1 net1 CLKIN sky130_fd_pr__cap_mim_m3_1 W=3e+07u L=3e+07u MF=100 m=100
XC2 VOUT GND sky130_fd_pr__cap_mim_m3_1 W=3e+07u L=3e+07u MF=100 m=100
.ends

.GLOBAL GND
** flattened .save nodes
.end
