magic
tech sky130A
timestamp 1635946216
<< error_p >>
rect -10 519 -9 536
rect 8 519 10 536
rect -73 467 -56 468
rect 56 467 73 468
rect -73 459 -56 460
rect 56 459 73 460
rect -73 440 -56 441
rect 56 440 73 441
rect -73 433 -56 434
rect 56 433 73 434
rect -73 423 -56 424
rect 56 423 73 424
rect -73 404 -56 405
rect 56 404 73 405
rect -73 399 -56 400
rect 56 399 73 400
rect -73 387 -56 388
rect 56 387 73 388
rect -73 368 -56 369
rect 56 368 73 369
rect -73 365 -56 366
rect 56 365 73 366
rect -73 351 -56 352
rect 56 351 73 352
rect -73 331 -56 333
rect 56 331 73 333
rect -73 315 -56 316
rect 56 315 73 316
rect -73 296 -56 298
rect 56 296 73 298
rect -73 279 -56 280
rect 56 279 73 280
rect -73 263 -56 264
rect 56 263 73 264
rect -73 260 -56 261
rect 56 260 73 261
rect -73 243 -56 244
rect 56 243 73 244
rect -73 229 -56 230
rect 56 229 73 230
rect -73 224 -56 225
rect 56 224 73 225
rect -73 207 -56 208
rect 56 207 73 208
rect -73 195 -56 196
rect 56 195 73 196
rect -73 188 -56 189
rect 56 188 73 189
rect -73 171 -56 172
rect 56 171 73 172
rect -73 161 -56 162
rect 56 161 73 162
rect -73 152 -56 153
rect 56 152 73 153
rect -73 135 -56 136
rect 56 135 73 136
rect -73 127 -56 128
rect 56 127 73 128
rect -73 116 -56 117
rect 56 116 73 117
rect -73 99 -56 100
rect 56 99 73 100
rect -73 93 -56 94
rect 56 93 73 94
rect -73 80 -56 81
rect 56 80 73 81
rect -73 63 -56 64
rect 56 63 73 64
rect -73 59 -56 60
rect 56 59 73 60
rect -73 44 -56 45
rect 56 44 73 45
rect -73 27 -56 28
rect 56 27 73 28
rect -73 25 -56 26
rect 56 25 73 26
rect -73 8 -56 9
rect 56 8 73 9
rect -73 -9 -56 -8
rect 56 -9 73 -8
rect -73 -28 -56 -27
rect 56 -28 73 -27
rect -73 -43 -56 -42
rect 56 -43 73 -42
rect -73 -45 -56 -44
rect 56 -45 73 -44
rect -73 -64 -56 -63
rect 56 -64 73 -63
rect -73 -77 -56 -76
rect 56 -77 73 -76
rect -73 -81 -56 -80
rect 56 -81 73 -80
rect -73 -100 -56 -99
rect 56 -100 73 -99
rect -73 -111 -56 -110
rect 56 -111 73 -110
rect -73 -117 -56 -116
rect 56 -117 73 -116
rect -73 -136 -56 -135
rect 56 -136 73 -135
rect -73 -145 -56 -144
rect 56 -145 73 -144
rect -73 -153 -56 -152
rect 56 -153 73 -152
rect -73 -172 -56 -171
rect 56 -172 73 -171
rect -73 -179 -56 -178
rect 56 -179 73 -178
rect -73 -189 -56 -188
rect 56 -189 73 -188
rect -73 -208 -56 -207
rect 56 -208 73 -207
rect -73 -213 -56 -212
rect 56 -213 73 -212
rect -73 -225 -56 -224
rect 56 -225 73 -224
rect -73 -244 -56 -243
rect 56 -244 73 -243
rect -73 -247 -56 -246
rect 56 -247 73 -246
rect -73 -261 -56 -260
rect 56 -261 73 -260
rect -73 -281 -56 -279
rect 56 -281 73 -279
rect -73 -297 -56 -296
rect 56 -297 73 -296
rect -73 -316 -56 -314
rect 56 -316 73 -314
rect -73 -333 -56 -332
rect 56 -333 73 -332
rect -73 -349 -56 -348
rect 56 -349 73 -348
rect -73 -352 -56 -351
rect 56 -352 73 -351
rect -73 -369 -56 -368
rect 56 -369 73 -368
rect -73 -383 -56 -382
rect 56 -383 73 -382
rect -73 -388 -56 -387
rect 56 -388 73 -387
rect -73 -405 -56 -404
rect 56 -405 73 -404
rect -73 -417 -56 -416
rect 56 -417 73 -416
rect -73 -424 -56 -423
rect 56 -424 73 -423
rect -73 -441 -56 -440
rect 56 -441 73 -440
rect -73 -451 -56 -450
rect 56 -451 73 -450
rect -73 -460 -56 -459
rect 56 -460 73 -459
rect -10 -536 -9 -519
rect 8 -536 10 -519
<< pwell >>
rect -92 -513 92 513
<< mvnmos >>
rect -50 -500 50 500
<< mvndiff >>
rect -79 485 -50 500
rect -79 467 -73 485
rect -56 467 -50 485
rect -79 451 -50 467
rect -79 433 -73 451
rect -56 433 -50 451
rect -79 417 -50 433
rect -79 399 -73 417
rect -56 399 -50 417
rect -79 383 -50 399
rect -79 365 -73 383
rect -56 365 -50 383
rect -79 349 -50 365
rect -79 331 -73 349
rect -56 331 -50 349
rect -79 315 -50 331
rect -79 297 -73 315
rect -56 297 -50 315
rect -79 281 -50 297
rect -79 263 -73 281
rect -56 263 -50 281
rect -79 247 -50 263
rect -79 229 -73 247
rect -56 229 -50 247
rect -79 213 -50 229
rect -79 195 -73 213
rect -56 195 -50 213
rect -79 179 -50 195
rect -79 161 -73 179
rect -56 161 -50 179
rect -79 145 -50 161
rect -79 127 -73 145
rect -56 127 -50 145
rect -79 111 -50 127
rect -79 93 -73 111
rect -56 93 -50 111
rect -79 77 -50 93
rect -79 59 -73 77
rect -56 59 -50 77
rect -79 43 -50 59
rect -79 25 -73 43
rect -56 25 -50 43
rect -79 9 -50 25
rect -79 -9 -73 9
rect -56 -9 -50 9
rect -79 -25 -50 -9
rect -79 -43 -73 -25
rect -56 -43 -50 -25
rect -79 -59 -50 -43
rect -79 -77 -73 -59
rect -56 -77 -50 -59
rect -79 -93 -50 -77
rect -79 -111 -73 -93
rect -56 -111 -50 -93
rect -79 -127 -50 -111
rect -79 -145 -73 -127
rect -56 -145 -50 -127
rect -79 -161 -50 -145
rect -79 -179 -73 -161
rect -56 -179 -50 -161
rect -79 -195 -50 -179
rect -79 -213 -73 -195
rect -56 -213 -50 -195
rect -79 -229 -50 -213
rect -79 -247 -73 -229
rect -56 -247 -50 -229
rect -79 -263 -50 -247
rect -79 -281 -73 -263
rect -56 -281 -50 -263
rect -79 -297 -50 -281
rect -79 -315 -73 -297
rect -56 -315 -50 -297
rect -79 -331 -50 -315
rect -79 -349 -73 -331
rect -56 -349 -50 -331
rect -79 -365 -50 -349
rect -79 -383 -73 -365
rect -56 -383 -50 -365
rect -79 -399 -50 -383
rect -79 -417 -73 -399
rect -56 -417 -50 -399
rect -79 -433 -50 -417
rect -79 -451 -73 -433
rect -56 -451 -50 -433
rect -79 -467 -50 -451
rect -79 -485 -73 -467
rect -56 -485 -50 -467
rect -79 -500 -50 -485
rect 50 485 79 500
rect 50 467 56 485
rect 73 467 79 485
rect 50 451 79 467
rect 50 433 56 451
rect 73 433 79 451
rect 50 417 79 433
rect 50 399 56 417
rect 73 399 79 417
rect 50 383 79 399
rect 50 365 56 383
rect 73 365 79 383
rect 50 349 79 365
rect 50 331 56 349
rect 73 331 79 349
rect 50 315 79 331
rect 50 297 56 315
rect 73 297 79 315
rect 50 281 79 297
rect 50 263 56 281
rect 73 263 79 281
rect 50 247 79 263
rect 50 229 56 247
rect 73 229 79 247
rect 50 213 79 229
rect 50 195 56 213
rect 73 195 79 213
rect 50 179 79 195
rect 50 161 56 179
rect 73 161 79 179
rect 50 145 79 161
rect 50 127 56 145
rect 73 127 79 145
rect 50 111 79 127
rect 50 93 56 111
rect 73 93 79 111
rect 50 77 79 93
rect 50 59 56 77
rect 73 59 79 77
rect 50 43 79 59
rect 50 25 56 43
rect 73 25 79 43
rect 50 9 79 25
rect 50 -9 56 9
rect 73 -9 79 9
rect 50 -25 79 -9
rect 50 -43 56 -25
rect 73 -43 79 -25
rect 50 -59 79 -43
rect 50 -77 56 -59
rect 73 -77 79 -59
rect 50 -93 79 -77
rect 50 -111 56 -93
rect 73 -111 79 -93
rect 50 -127 79 -111
rect 50 -145 56 -127
rect 73 -145 79 -127
rect 50 -161 79 -145
rect 50 -179 56 -161
rect 73 -179 79 -161
rect 50 -195 79 -179
rect 50 -213 56 -195
rect 73 -213 79 -195
rect 50 -229 79 -213
rect 50 -247 56 -229
rect 73 -247 79 -229
rect 50 -263 79 -247
rect 50 -281 56 -263
rect 73 -281 79 -263
rect 50 -297 79 -281
rect 50 -315 56 -297
rect 73 -315 79 -297
rect 50 -331 79 -315
rect 50 -349 56 -331
rect 73 -349 79 -331
rect 50 -365 79 -349
rect 50 -383 56 -365
rect 73 -383 79 -365
rect 50 -399 79 -383
rect 50 -417 56 -399
rect 73 -417 79 -399
rect 50 -433 79 -417
rect 50 -451 56 -433
rect 73 -451 79 -433
rect 50 -467 79 -451
rect 50 -485 56 -467
rect 73 -485 79 -467
rect 50 -500 79 -485
<< mvndiffc >>
rect -73 467 -56 485
rect -73 433 -56 451
rect -73 399 -56 417
rect -73 365 -56 383
rect -73 331 -56 349
rect -73 297 -56 315
rect -73 263 -56 281
rect -73 229 -56 247
rect -73 195 -56 213
rect -73 161 -56 179
rect -73 127 -56 145
rect -73 93 -56 111
rect -73 59 -56 77
rect -73 25 -56 43
rect -73 -9 -56 9
rect -73 -43 -56 -25
rect -73 -77 -56 -59
rect -73 -111 -56 -93
rect -73 -145 -56 -127
rect -73 -179 -56 -161
rect -73 -213 -56 -195
rect -73 -247 -56 -229
rect -73 -281 -56 -263
rect -73 -315 -56 -297
rect -73 -349 -56 -331
rect -73 -383 -56 -365
rect -73 -417 -56 -399
rect -73 -451 -56 -433
rect -73 -485 -56 -467
rect 56 467 73 485
rect 56 433 73 451
rect 56 399 73 417
rect 56 365 73 383
rect 56 331 73 349
rect 56 297 73 315
rect 56 263 73 281
rect 56 229 73 247
rect 56 195 73 213
rect 56 161 73 179
rect 56 127 73 145
rect 56 93 73 111
rect 56 59 73 77
rect 56 25 73 43
rect 56 -9 73 9
rect 56 -43 73 -25
rect 56 -77 73 -59
rect 56 -111 73 -93
rect 56 -145 73 -127
rect 56 -179 73 -161
rect 56 -213 73 -195
rect 56 -247 73 -229
rect 56 -281 73 -263
rect 56 -315 73 -297
rect 56 -349 73 -331
rect 56 -383 73 -365
rect 56 -417 73 -399
rect 56 -451 73 -433
rect 56 -485 73 -467
<< poly >>
rect -50 536 50 544
rect -50 519 -26 536
rect -8 519 8 536
rect 26 519 50 536
rect -50 500 50 519
rect -50 -519 50 -500
rect -50 -536 -26 -519
rect -8 -536 8 -519
rect 26 -536 50 -519
rect -50 -544 50 -536
<< polycont >>
rect -26 519 -8 536
rect 8 519 26 536
rect -26 -536 -8 -519
rect 8 -536 26 -519
<< locali >>
rect -50 519 -27 536
rect -8 519 8 536
rect 27 519 50 536
rect -73 485 -56 502
rect -73 451 -56 459
rect -73 417 -56 423
rect -73 383 -56 387
rect -73 349 -56 351
rect -73 261 -56 263
rect -73 225 -56 229
rect -73 189 -56 195
rect -73 153 -56 161
rect -73 117 -56 127
rect -73 81 -56 93
rect -73 45 -56 59
rect -73 9 -56 25
rect -73 -25 -56 -9
rect -73 -59 -56 -45
rect -73 -93 -56 -81
rect -73 -127 -56 -117
rect -73 -161 -56 -153
rect -73 -195 -56 -189
rect -73 -229 -56 -225
rect -73 -263 -56 -261
rect -73 -351 -56 -349
rect -73 -387 -56 -383
rect -73 -423 -56 -417
rect -73 -459 -56 -451
rect -73 -502 -56 -485
rect 56 485 73 502
rect 56 451 73 459
rect 56 417 73 423
rect 56 383 73 387
rect 56 349 73 351
rect 56 261 73 263
rect 56 225 73 229
rect 56 189 73 195
rect 56 153 73 161
rect 56 117 73 127
rect 56 81 73 93
rect 56 45 73 59
rect 56 9 73 25
rect 56 -25 73 -9
rect 56 -59 73 -45
rect 56 -93 73 -81
rect 56 -127 73 -117
rect 56 -161 73 -153
rect 56 -195 73 -189
rect 56 -229 73 -225
rect 56 -263 73 -261
rect 56 -351 73 -349
rect 56 -387 73 -383
rect 56 -423 73 -417
rect 56 -459 73 -451
rect 56 -502 73 -485
rect -50 -536 -27 -519
rect -8 -536 8 -519
rect 27 -536 50 -519
<< viali >>
rect -27 519 -26 536
rect -26 519 -9 536
rect 9 519 26 536
rect 26 519 27 536
rect -73 467 -56 477
rect -73 459 -56 467
rect -73 433 -56 441
rect -73 423 -56 433
rect -73 399 -56 405
rect -73 387 -56 399
rect -73 365 -56 369
rect -73 351 -56 365
rect -73 331 -56 333
rect -73 315 -56 331
rect -73 281 -56 297
rect -73 279 -56 281
rect -73 247 -56 261
rect -73 243 -56 247
rect -73 213 -56 225
rect -73 207 -56 213
rect -73 179 -56 189
rect -73 171 -56 179
rect -73 145 -56 153
rect -73 135 -56 145
rect -73 111 -56 117
rect -73 99 -56 111
rect -73 77 -56 81
rect -73 63 -56 77
rect -73 43 -56 45
rect -73 27 -56 43
rect -73 -9 -56 9
rect -73 -43 -56 -27
rect -73 -45 -56 -43
rect -73 -77 -56 -63
rect -73 -81 -56 -77
rect -73 -111 -56 -99
rect -73 -117 -56 -111
rect -73 -145 -56 -135
rect -73 -153 -56 -145
rect -73 -179 -56 -171
rect -73 -189 -56 -179
rect -73 -213 -56 -207
rect -73 -225 -56 -213
rect -73 -247 -56 -243
rect -73 -261 -56 -247
rect -73 -281 -56 -279
rect -73 -297 -56 -281
rect -73 -331 -56 -315
rect -73 -333 -56 -331
rect -73 -365 -56 -351
rect -73 -369 -56 -365
rect -73 -399 -56 -387
rect -73 -405 -56 -399
rect -73 -433 -56 -423
rect -73 -441 -56 -433
rect -73 -467 -56 -459
rect -73 -477 -56 -467
rect 56 467 73 477
rect 56 459 73 467
rect 56 433 73 441
rect 56 423 73 433
rect 56 399 73 405
rect 56 387 73 399
rect 56 365 73 369
rect 56 351 73 365
rect 56 331 73 333
rect 56 315 73 331
rect 56 281 73 297
rect 56 279 73 281
rect 56 247 73 261
rect 56 243 73 247
rect 56 213 73 225
rect 56 207 73 213
rect 56 179 73 189
rect 56 171 73 179
rect 56 145 73 153
rect 56 135 73 145
rect 56 111 73 117
rect 56 99 73 111
rect 56 77 73 81
rect 56 63 73 77
rect 56 43 73 45
rect 56 27 73 43
rect 56 -9 73 9
rect 56 -43 73 -27
rect 56 -45 73 -43
rect 56 -77 73 -63
rect 56 -81 73 -77
rect 56 -111 73 -99
rect 56 -117 73 -111
rect 56 -145 73 -135
rect 56 -153 73 -145
rect 56 -179 73 -171
rect 56 -189 73 -179
rect 56 -213 73 -207
rect 56 -225 73 -213
rect 56 -247 73 -243
rect 56 -261 73 -247
rect 56 -281 73 -279
rect 56 -297 73 -281
rect 56 -331 73 -315
rect 56 -333 73 -331
rect 56 -365 73 -351
rect 56 -369 73 -365
rect 56 -399 73 -387
rect 56 -405 73 -399
rect 56 -433 73 -423
rect 56 -441 73 -433
rect 56 -467 73 -459
rect 56 -477 73 -467
rect -27 -536 -26 -519
rect -26 -536 -9 -519
rect 9 -536 26 -519
rect 26 -536 27 -519
<< metal1 >>
rect -48 536 48 539
rect -48 519 -27 536
rect -9 519 9 536
rect 27 519 48 536
rect -48 516 48 519
rect -76 477 -53 500
rect -76 459 -73 477
rect -56 459 -53 477
rect -76 441 -53 459
rect -76 423 -73 441
rect -56 423 -53 441
rect -76 405 -53 423
rect -76 387 -73 405
rect -56 387 -53 405
rect -76 369 -53 387
rect -76 351 -73 369
rect -56 351 -53 369
rect -76 333 -53 351
rect -76 315 -73 333
rect -56 315 -53 333
rect -76 297 -53 315
rect -76 279 -73 297
rect -56 279 -53 297
rect -76 261 -53 279
rect -76 243 -73 261
rect -56 243 -53 261
rect -76 225 -53 243
rect -76 207 -73 225
rect -56 207 -53 225
rect -76 189 -53 207
rect -76 171 -73 189
rect -56 171 -53 189
rect -76 153 -53 171
rect -76 135 -73 153
rect -56 135 -53 153
rect -76 117 -53 135
rect -76 99 -73 117
rect -56 99 -53 117
rect -76 81 -53 99
rect -76 63 -73 81
rect -56 63 -53 81
rect -76 45 -53 63
rect -76 27 -73 45
rect -56 27 -53 45
rect -76 9 -53 27
rect -76 -9 -73 9
rect -56 -9 -53 9
rect -76 -27 -53 -9
rect -76 -45 -73 -27
rect -56 -45 -53 -27
rect -76 -63 -53 -45
rect -76 -81 -73 -63
rect -56 -81 -53 -63
rect -76 -99 -53 -81
rect -76 -117 -73 -99
rect -56 -117 -53 -99
rect -76 -135 -53 -117
rect -76 -153 -73 -135
rect -56 -153 -53 -135
rect -76 -171 -53 -153
rect -76 -189 -73 -171
rect -56 -189 -53 -171
rect -76 -207 -53 -189
rect -76 -225 -73 -207
rect -56 -225 -53 -207
rect -76 -243 -53 -225
rect -76 -261 -73 -243
rect -56 -261 -53 -243
rect -76 -279 -53 -261
rect -76 -297 -73 -279
rect -56 -297 -53 -279
rect -76 -315 -53 -297
rect -76 -333 -73 -315
rect -56 -333 -53 -315
rect -76 -351 -53 -333
rect -76 -369 -73 -351
rect -56 -369 -53 -351
rect -76 -387 -53 -369
rect -76 -405 -73 -387
rect -56 -405 -53 -387
rect -76 -423 -53 -405
rect -76 -441 -73 -423
rect -56 -441 -53 -423
rect -76 -459 -53 -441
rect -76 -477 -73 -459
rect -56 -477 -53 -459
rect -76 -500 -53 -477
rect 53 477 76 500
rect 53 459 56 477
rect 73 459 76 477
rect 53 441 76 459
rect 53 423 56 441
rect 73 423 76 441
rect 53 405 76 423
rect 53 387 56 405
rect 73 387 76 405
rect 53 369 76 387
rect 53 351 56 369
rect 73 351 76 369
rect 53 333 76 351
rect 53 315 56 333
rect 73 315 76 333
rect 53 297 76 315
rect 53 279 56 297
rect 73 279 76 297
rect 53 261 76 279
rect 53 243 56 261
rect 73 243 76 261
rect 53 225 76 243
rect 53 207 56 225
rect 73 207 76 225
rect 53 189 76 207
rect 53 171 56 189
rect 73 171 76 189
rect 53 153 76 171
rect 53 135 56 153
rect 73 135 76 153
rect 53 117 76 135
rect 53 99 56 117
rect 73 99 76 117
rect 53 81 76 99
rect 53 63 56 81
rect 73 63 76 81
rect 53 45 76 63
rect 53 27 56 45
rect 73 27 76 45
rect 53 9 76 27
rect 53 -9 56 9
rect 73 -9 76 9
rect 53 -27 76 -9
rect 53 -45 56 -27
rect 73 -45 76 -27
rect 53 -63 76 -45
rect 53 -81 56 -63
rect 73 -81 76 -63
rect 53 -99 76 -81
rect 53 -117 56 -99
rect 73 -117 76 -99
rect 53 -135 76 -117
rect 53 -153 56 -135
rect 73 -153 76 -135
rect 53 -171 76 -153
rect 53 -189 56 -171
rect 73 -189 76 -171
rect 53 -207 76 -189
rect 53 -225 56 -207
rect 73 -225 76 -207
rect 53 -243 76 -225
rect 53 -261 56 -243
rect 73 -261 76 -243
rect 53 -279 76 -261
rect 53 -297 56 -279
rect 73 -297 76 -279
rect 53 -315 76 -297
rect 53 -333 56 -315
rect 73 -333 76 -315
rect 53 -351 76 -333
rect 53 -369 56 -351
rect 73 -369 76 -351
rect 53 -387 76 -369
rect 53 -405 56 -387
rect 73 -405 76 -387
rect 53 -423 76 -405
rect 53 -441 56 -423
rect 73 -441 76 -423
rect 53 -459 76 -441
rect 53 -477 56 -459
rect 73 -477 76 -459
rect 53 -500 76 -477
rect -48 -519 48 -516
rect -48 -536 -27 -519
rect -9 -536 9 -519
rect 27 -536 48 -519
rect -48 -539 48 -536
<< end >>
