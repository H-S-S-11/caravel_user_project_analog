  X �    ' �    '  LIB  >A�7KƧ�9D�/��ZX �    ' �    '  contact$2     B  , ,������������   U����   U����������������      B  , ,   _����   _   U  	   U  	����   _����      C   ,�������[����   �  Y   �  Y���[�������[      A  , ,������3���   �  �   �  ����3������3     �    ' �    '  (sky130_fd_pr__nfet_g5v0d10v5_9A4VCP     D   ,���   (���     �    �  (���   (      D   ,������x���  �����  ��������x������x      D   ,  ���x    �  �  �  ����x  ���x      D   ,��� ������� ����  �����  �������� ����      B  , ,���  F���  �����  �����  F���  F      B  , ,   U  F   U  �   �  �   �  F   U  F      B  , ,���&  C���&  �����  �����  C���&  C      B  , ,  0  C  0  �  �  �  �  C  0  C      B  , ,���&  ����&  �����  �����  ����&  �      B  , ,  0  �  0  �  �  �  �  �  0  �      B  , ,���&  ����&  E����  E����  ����&  �      B  , ,  0  �  0  E  �  E  �  �  0  �      B  , ,���&  G���&  �����  �����  G���&  G      B  , ,  0  G  0  �  �  �  �  G  0  G      B  , ,���&  ����&  �����  �����  ����&  �      B  , ,  0  �  0  �  �  �  �  �  0  �      B  , ,���&  ����&  I����  I����  ����&  �      B  , ,  0  �  0  I  �  I  �  �  0  �      B  , ,���&  
K���&  
�����  
�����  
K���&  
K      B  , ,  0  
K  0  
�  �  
�  �  
K  0  
K      B  , ,���&  ����&  	�����  	�����  ����&  �      B  , ,  0  �  0  	�  �  	�  �  �  0  �      B  , ,���&  ����&  M����  M����  ����&  �      B  , ,  0  �  0  M  �  M  �  �  0  �      B  , ,���&  O���&  �����  �����  O���&  O      B  , ,  0  O  0  �  �  �  �  O  0  O      B  , ,���&  ����&  �����  �����  ����&  �      B  , ,  0  �  0  �  �  �  �  �  0  �      B  , ,���&  ����&  Q����  Q����  ����&  �      B  , ,  0  �  0  Q  �  Q  �  �  0  �      B  , ,���&  S���&  �����  �����  S���&  S      B  , ,  0  S  0  �  �  �  �  S  0  S      B  , ,���&   ����&  �����  �����   ����&   �      B  , ,  0   �  0  �  �  �  �   �  0   �      B  , ,���&�������&   U����   U�����������&����      B  , ,  0����  0   U  �   U  �����  0����      B  , ,���&���W���&�����������������W���&���W      B  , ,  0���W  0���  ����  ����W  0���W      B  , ,���&������&����������������������&���      B  , ,  0���  0����  �����  ����  0���      B  , ,���&�������&���Y�������Y�����������&����      B  , ,  0����  0���Y  ����Y  �����  0����      B  , ,���&���[���&�����������������[���&���[      B  , ,  0���[  0���  ����  ����[  0���[      B  , ,���&������&����������������������&���      B  , ,  0���  0����  �����  ����  0���      B  , ,���&�������&���]�������]�����������&����      B  , ,  0����  0���]  ����]  �����  0����      B  , ,���&���_���&���	�������	�������_���&���_      B  , ,  0���_  0���	  ����	  ����_  0���_      B  , ,���&������&����������������������&���      B  , ,  0���  0����  �����  ����  0���      B  , ,���&������&���a�������a����������&���      B  , ,  0���  0���a  ����a  ����  0���      B  , ,���&���c���&�����������������c���&���c      B  , ,  0���c  0���  ����  ����c  0���c      B  , ,���&������&��������������������&���      B  , ,  0���  0���  ����  ����  0���      B  , ,���&������&���e�������e����������&���      B  , ,  0���  0���e  ����e  ����  0���      B  , ,���&���g���&�����������������g���&���g      B  , ,  0���g  0���  ����  ����g  0���g      B  , ,���&������&��������������������&���      B  , ,  0���  0���  ����  ����  0���      B  , ,��������������������������������      B  , ,   U���   U���   ����   ����   U���      C   ,���  F���  �  �  �  �  F���  F      C   ,���&���d���&  �����  ��������d���&���d      C   ,  0���d  0  �  �  �  ����d  0���d      C   ,������������  ����  ����������      C  , ,����  F����  �����  �����  F����  F      C  , ,   _  F   _  �  	  �  	  F   _  F      C  , ,���&  ����&  �����  �����  ����&  �      C  , ,  0  �  0  �  �  �  �  �  0  �      C  , ,���&  ����&  5����  5����  ����&  �      C  , ,  0  �  0  5  �  5  �  �  0  �      C  , ,���&  #���&  �����  �����  #���&  #      C  , ,  0  #  0  �  �  �  �  #  0  #      C  , ,���&  ����&  e����  e����  ����&  �      C  , ,  0  �  0  e  �  e  �  �  0  �      C  , ,���&  S���&  �����  �����  S���&  S      C  , ,  0  S  0  �  �  �  �  S  0  S      C  , ,���&  
����&  �����  �����  
����&  
�      C  , ,  0  
�  0  �  �  �  �  
�  0  
�      C  , ,���&  	����&  
-����  
-����  	����&  	�      C  , ,  0  	�  0  
-  �  
-  �  	�  0  	�      C  , ,���&  ���&  �����  �����  ���&        C  , ,  0    0  �  �  �  �    0        C  , ,���&  ����&  ]����  ]����  ����&  �      C  , ,  0  �  0  ]  �  ]  �  �  0  �      C  , ,���&  K���&  �����  �����  K���&  K      C  , ,  0  K  0  �  �  �  �  K  0  K      C  , ,���&  ����&  �����  �����  ����&  �      C  , ,  0  �  0  �  �  �  �  �  0  �      C  , ,���&  {���&  %����  %����  {���&  {      C  , ,  0  {  0  %  �  %  �  {  0  {      C  , ,���&  ���&  �����  �����  ���&        C  , ,  0    0  �  �  �  �    0        C  , ,���&�������&   U����   U�����������&����      C  , ,  0����  0   U  �   U  �����  0����      C  , ,���&���C���&�������������������C���&���C      C  , ,  0���C  0����  �����  ����C  0���C      C  , ,���&�������&�����������������������&����      C  , ,  0����  0����  �����  �����  0����      C  , ,���&���s���&�����������������s���&���s      C  , ,  0���s  0���  ����  ����s  0���s      C  , ,���&������&����������������������&���      C  , ,  0���  0����  �����  ����  0���      C  , ,���&�������&���M�������M�����������&����      C  , ,  0����  0���M  ����M  �����  0����      C  , ,���&���;���&�������������������;���&���;      C  , ,  0���;  0����  �����  ����;  0���;      C  , ,���&�������&���}�������}�����������&����      C  , ,  0����  0���}  ����}  �����  0����      C  , ,���&���k���&�����������������k���&���k      C  , ,  0���k  0���  ����  ����k  0���k      C  , ,���&������&��������������������&���      C  , ,  0���  0���  ����  ����  0���      C  , ,���&������&���E�������E����������&���      C  , ,  0���  0���E  ����E  ����  0���      C  , ,���&���3���&�������������������3���&���3      C  , ,  0���3  0����  �����  ����3  0���3      C  , ,���&�������&���u�������u�����������&����      C  , ,  0����  0���u  ����u  �����  0����      C  , ,���&���c���&�����������������c���&���c      C  , ,  0���c  0���  ����  ����c  0���c      C  , ,�����������������������������������      C  , ,   _���   _���  	���  	���   _���      A   ,�������x����  �    �  ���x�������x      B   ,����������  @  �  @  ������������      K   ,���1������1  A  �  A  �������1���      _   ,����  �����  T  c  T  c  �����  �      _   ,��������������  c���  c����������      ]  , ,���m�������m    �    ��������m����      }   ,���1������1  A  �  A  �������1���     �    ' �    '  contact$4     D   ,�������`����   �  @   �  @���`�������`      D  , ,����������   K����   K���������������      D  , ,   U����   U   K   �   K   �����   U����      E   ,�������`����   �  @   �  @���`�������`     �    ' �    '  (sky130_fd_pr__pfet_g5v0d10v5_QSRSHK     D   ,���,  ����,  �  �  �  �  ����,  �      D   ,���������  �����  ��������������      D   ,  ���    �  �  �  ����  ���      D   ,���,���e���,���K  ����K  ����e���,���e      B  , ,���  ����  }����  }����  ����  �      B  , ,���W  ����W  }���  }���  ����W  �      B  , ,����  �����  }   U  }   U  �����  �      B  , ,   �  �   �  }  �  }  �  �   �  �      B  , ,  S  �  S  }  �  }  �  �  S  �      B  , ,���2  ����2  �����  �����  ����2  �      B  , ,  $  �  $  �  �  �  �  �  $  �      B  , ,���2  ����2  S����  S����  ����2  �      B  , ,  $  �  $  S  �  S  �  �  $  �      B  , ,���2   U���2   �����   �����   U���2   U      B  , ,  $   U  $   �  �   �  �   U  $   U      B  , ,���2������2����������������������2���      B  , ,  $���  $����  �����  ����  $���      B  , ,���2�������2���W�������W�����������2����      B  , ,  $����  $���W  ����W  �����  $����      B  , ,���2���Y���2�����������������Y���2���Y      B  , ,  $���Y  $���  ����  ����Y  $���Y      B  , ,�������������-�������-���������������      B  , ,���W�������W���-������-����������W����      B  , ,���������������-   U���-   U������������      B  , ,   �����   ����-  ����-  �����   �����      B  , ,  S����  S���-  ����-  �����  S����      C   ,���  ����  }  �  }  �  ����  �      C   ,���2������2  �����  �����������2���      C   ,  $���  $  �  �  �  ����  $���      C   ,�������������-  ����-  ������������      C  , ,����  �����  }����  }����  �����  �      C  , ,���C  ����C  }����  }����  ����C  �      C  , ,����  �����  }   U  }   U  �����  �      C  , ,    �    }  �  }  �  �    �      C  , ,  {  �  {  }  %  }  %  �  {  �      C  , ,���2  {���2  %����  %����  {���2  {      C  , ,  $  {  $  %  �  %  �  {  $  {      C  , ,���2  ���2  �����  �����  ���2        C  , ,  $    $  �  �  �  �    $        C  , ,���2�������2   U����   U�����������2����      C  , ,  $����  $   U  �   U  �����  $����      C  , ,���2���C���2�������������������C���2���C      C  , ,  $���C  $����  �����  ����C  $���C      C  , ,���2�������2�����������������������2����      C  , ,  $����  $����  �����  �����  $����      C  , ,���������������-�������-����������������      C  , ,���C�������C���-�������-�����������C����      C  , ,���������������-   U���-   U������������      C  , ,  ����  ���-  ����-  �����  ����      C  , ,  {����  {���-  %���-  %����  {����      A   ,�����������  �  
  �  
����������      B   ,������3���  �  �  �  ����3������3      K   ,���B  ����B  �  �  �  �  ����B  �      K   ,���=���_���=  �  �  �  ����_���=���_      K   ,���B���$���B���_  ����_  ����$���B���$      _   ,����  o����  �  a  �  a  o����  o      _   ,���������������  a����  a����������      ^   ,���y�������y  e  �  e  ��������y����      @   ,���B�������B  
n  �  
n  ��������B����     �    ' �    '  (sky130_fd_pr__nfet_g5v0d10v5_DPU6YB     D   ,���,  ����,  z  �  z  �  ����,  �      D   ,���������  �����  ��������������      D   ,  ���    �  �  �  ����  ���      D   ,���,�������,���l  ����l  ��������,����      B  , ,���  ����  \����  \����  ����  �      B  , ,���W  ����W  \���  \���  ����W  �      B  , ,����  �����  \   U  \   U  �����  �      B  , ,   �  �   �  \  �  \  �  �   �  �      B  , ,  S  �  S  \  �  \  �  �  S  �      B  , ,���2   ����2  �����  �����   ����2   �      B  , ,  $   �  $  �  �  �  �   �  $   �      B  , ,���2�������2   U����   U�����������2����      B  , ,  $����  $   U  �   U  �����  $����      B  , ,���2���W���2�����������������W���2���W      B  , ,  $���W  $���  ����  ����W  $���W      B  , ,�������������N�������N���������������      B  , ,���W�������W���N������N����������W����      B  , ,���������������N   U���N   U������������      B  , ,   �����   ����N  ����N  �����   �����      B  , ,  S����  S���N  ����N  �����  S����      C   ,���  ����  \  �  \  �  ����  �      C   ,���2�������2  ����  �����������2����      C   ,  $����  $    �    �����  $����      C   ,�������������N  ����N  ������������      C  , ,����  �����  \����  \����  �����  �      C  , ,���C  ����C  \����  \����  ����C  �      C  , ,����  �����  \   U  \   U  �����  �      C  , ,    �    \  �  \  �  �    �      C  , ,  {  �  {  \  %  \  %  �  {  �      C  , ,���2   _���2  	����  	����   _���2   _      C  , ,  $   _  $  	  �  	  �   _  $   _      C  , ,���2�������2�����������������������2����      C  , ,  $����  $����  �����  �����  $����      C  , ,���������������N�������N����������������      C  , ,���C�������C���N�������N�����������C����      C  , ,���������������N   U���N   U������������      C  , ,  ����  ���N  ����N  �����  ����      C  , ,  {����  {���N  %���N  %����  {����      A   ,�����������  �  
  �  
����������      B   ,������T���  �  �  �  ����T������T      K   ,���=���S���=  �  �  �  ����S���=���S      _   ,����  N����  �  a  �  a  N����  N      _   ,�������@��������  a����  a���@�������@      ]  , ,���y�������y  q  �  q  ��������y����      }   ,���=���S���=  �  �  �  ����S���=���S     �    ' �    '  contact$3     D   ,�������o����   �  E   �  E���o�������o      C   ,�������[����   �  Y   �  Y���[�������[      C  , ,������������   U����   U����������������      C  , ,   _����   _   U  	   U  	����   _����     �    ' �    '  nfet_w10_l1  
  (sky130_fd_pr__nfet_g5v0d10v5_9A4VCP  ����  �   
  contact$2  ����  (x   
  contact$4  ��������      D   ,��ͺ���<��ͺ  #
���b  #
���b���<��ͺ���<      D   ,���"�������"  -�����  -������������"����      D   ,���������������t��̢���t��̢������������      ^   ,��ȡ  &���ȡ  *!���G  *!���G  &���ȡ  &�     �    ' �    '  m2_pfet_w2_l2  
  contact$2  �������w   
  contact$3  �������w   
  contact$2  ����  �   
  contact$3  ����  �     (sky130_fd_pr__pfet_g5v0d10v5_QSRSHK                           �      D   ,���,  ����,  �  �  �  �  ����,  �      D   ,���{���s���{  ����  �������s���{���s      D   ,  ����!  �  �  �  �  ����!  ����!      D   ,������s������{  |���{  |���s������s      D   ,���  ����  �  |  �  |  ����  �      ]  , ,���������������  �����  �����������      ]  , ,����  w����  )  �  )  �  w����  w     �    ' �    '  contact    �    ' �    '  m2_nfet_w1_l2    contact$2     �������`�������`�������`     contact$3     �������`�������`�������`     contact$2     ����  �����  �����  �     contact$3     ����  �����  �����  �     (sky130_fd_pr__nfet_g5v0d10v5_DPU6YB     ��������������������  x      D   ,���I���)���I  ����  �������)���I���)      D   ,����������������������������������������      D   ,����  
�����  ����  ����  
�����  
�      D   ,�������j����  :���z  :���z���j�������j      D   ,�����������  
i    
i  ����������      ^   ,�������������������������������������      ^   ,����  
<����  �����  �����  
<����  
<     �    ' �    '  m10_nfet_w10_l1    nfet_w10_l1   
    D  �  ��  �  D  �      D   ,���f  /����f  2�  J  2�  J  /����f  /�      D   ,��������������+  R����+  R�����������      E   ,��Й������Й���Z  N����Z  N�������Й����      E   ,���  )T���  +H  N�  +H  N�  )T���  )T     �    ' �    '  amp    m2_pfet_w2_l2     ���%���  X�������%���     contact$4     ���W  N  X�  N���W  N      D   ,���)  ���)  �  BE  �  BE  ���)        D   ,������������5  N����5  N����������      E   ,���  T���  H  H�  H  H�  T���  T     �    ' �    '  current_mirror   m2_pfet_w2_l2     ����  �  �  �����  �     contact$4     ���      ���        D   ,����  	Q����  �����  �����  	Q����  	Q      D   ,���  ����  !  q  !  q  ����  �      E   ,���  
A���  �  �  �  �  
A���  
A     �    ' �    '  bias_current_mirror    m2_nfet_w1_l2   
  �������X  �F���X�������X     contact$4   
  ������/  ����/������/   
  contact  ���L  	�      D   ,���p��ٽ���p��܍������܍������ٽ���p��ٽ      D   ,���J���?���J��ʁ  ����ʁ  �����?���J���?      D   ,��������������������������������������      D   ,���:���?���:�����������������?���:���?      D   ,  	����  	���e  ����e  �����  	����      D   ,  ����e  �����  ������  �����e  ����e      D   ,  �����  ����e  	���e  	����  �����      D   ,  0 ����  0 ���e  2����e  2�����  0 ����      D   ,  C�����  C����e  F���e  F����  C�����      D   ,  W0����  W0���e  Y����e  Y�����  W0����      D   ,  j�����  j����e  m)���e  m)����  j�����      D   ,  ~@����  ~@���e  �����e  ������  ~@����      D   ,  ������  �����e  �9���e  �9����  ������      D   ,  �P����  �P���e  �����e  ������  �P����      E   ,���R���]���R���  �5���  �5���]���R���]     �    ' �    '  diff_pair    m10_nfet_w10_l1     ���'   Z 4�   Z���'   Z     �    ' �    '  (UNNAMED)$1  
  (sky130_fd_pr__nfet_g5v0d10v5_9A4VCP      @     �    ' �    '  myopamp  
  bias_current_mirror    )r  Cl   
  amp     xU   
  current_mirror   7�  �   
  diff_pair  ���  H�   
  contact$4    �<  z�      D   ,  0\  }2  0\  ��  2�  ��  2�  }2  0\  }2      D   ,  C�  }-  C�  ��  F}  ��  F}  }-  C�  }-      D   ,  2�  .�  2�  9  4�  9  4�  .�  2�  .�      D   ,  �3  .�  �3  18  �a  18  �a  .�  �3  .�      D   ,  �  18  �  b�  �a  b�  �a  18  �  18      D   ,  P�  �g  P�  ��  �B  ��  �B  �g  P�  �g      D   ,  :  ��  :  �&  SR  �&  SR  ��  :  ��      D   ,  P�  ��  P�  ��  SR  ��  SR  ��  P�  ��      D   ,  �a  F�  �a  M�  �7  M�  �7  F�  �a  F�      D   ,  0p  9  0p  <(  N�  <(  N�  9  0p  9      D   ,  C�  x�  C�  }-  F}  }-  F}  x�  C�  x�      D   ,  'L  x�  'L  }A  3  }A  3  x�  'L  x�      E   ,  ��  y�  ��  {�  �6  {�  �6  y�  ��  y�      D   ,  ��  F�  ��  M�  �#  M�  �#  F�  ��  F�      D   ,  �  	�  �  �  �  �  �  	�  �  	�      D   ,  �  ,�  �  /  '  /  '  ,�  �  ,�      D   ,  K  ��  K  �!   �  �!   �  ��  K  ��      D       m  � vdd       D       ��  Je out       D       `  � vss       D       �  -� bias      E   ,  �x  B�  �x  D9  ��  D9  ��  B�  �x  B�      E   ,  "�  B|  "�  D4  %�  D4  %�  B|  "�  B|      E   ,���R  r=���R  t;  ,  t;  ,  r=���R  r=      E   ,  K  r=  K  t;  M�  t;  M�  r=  K  r=      E       $,  CN in_n      E       ��  CI in_p      E       Lw  sK vss       E     ����  sK vss      �    ' �    '  devices  
  (sky130_fd_pr__nfet_g5v0d10v5_DPU6YB    
  �     �    ' �    '  (UNNAMED)  
  (sky130_fd_pr__pfet_g5v0d10v5_QSRSHK    
  �      