VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO myopamp
  CLASS BLOCK ;
  FOREIGN myopamp ;
  ORIGIN 45.995 -2.475 ;
  SIZE 215.245 BY 83.640 ;
  PIN vss
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 105.405 37.400 105.735 38.095 ;
        RECT 6.345 10.420 7.035 10.750 ;
        RECT 11.345 10.420 12.035 10.750 ;
        RECT 16.345 10.420 17.035 10.750 ;
        RECT 21.345 10.420 22.035 10.750 ;
        RECT 26.345 10.420 27.035 10.750 ;
        RECT 31.345 10.420 32.035 10.750 ;
        RECT 36.345 10.420 37.035 10.750 ;
        RECT 41.345 10.420 42.035 10.750 ;
        RECT 46.345 10.420 47.035 10.750 ;
        RECT 51.345 10.420 52.035 10.750 ;
        RECT 5.440 8.560 5.610 9.600 ;
        RECT 10.440 8.560 10.610 9.600 ;
        RECT 15.440 8.560 15.610 9.600 ;
        RECT 20.440 8.560 20.610 9.600 ;
        RECT 25.440 8.560 25.610 9.600 ;
        RECT 30.440 8.560 30.610 9.600 ;
        RECT 35.440 8.560 35.610 9.600 ;
        RECT 40.440 8.560 40.610 9.600 ;
        RECT 45.440 8.560 45.610 9.600 ;
        RECT 50.440 8.560 50.610 9.600 ;
        RECT 5.440 6.060 5.610 7.100 ;
        RECT 10.440 6.060 10.610 7.100 ;
        RECT 15.440 6.060 15.610 7.100 ;
        RECT 20.440 6.060 20.610 7.100 ;
        RECT 25.440 6.060 25.610 7.100 ;
        RECT 30.440 6.060 30.610 7.100 ;
        RECT 35.440 6.060 35.610 7.100 ;
        RECT 40.440 6.060 40.610 7.100 ;
        RECT 45.440 6.060 45.610 7.100 ;
        RECT 50.440 6.060 50.610 7.100 ;
        RECT 6.340 4.735 7.030 5.065 ;
        RECT 11.340 4.735 12.030 5.065 ;
        RECT 16.340 4.735 17.030 5.065 ;
        RECT 21.340 4.735 22.030 5.065 ;
        RECT 26.340 4.735 27.030 5.065 ;
        RECT 31.340 4.735 32.030 5.065 ;
        RECT 36.340 4.735 37.030 5.065 ;
        RECT 41.340 4.735 42.030 5.065 ;
        RECT 46.340 4.735 47.030 5.065 ;
        RECT 51.340 4.735 52.030 5.065 ;
      LAYER met1 ;
        RECT -23.970 13.065 -23.445 29.765 ;
        RECT 105.365 29.265 105.775 38.135 ;
        RECT 6.365 10.710 7.015 10.730 ;
        RECT 11.365 10.710 12.015 10.730 ;
        RECT 16.365 10.710 17.015 10.730 ;
        RECT 21.365 10.710 22.015 10.730 ;
        RECT 26.365 10.710 27.015 10.730 ;
        RECT 31.365 10.710 32.015 10.730 ;
        RECT 36.365 10.710 37.015 10.730 ;
        RECT 41.365 10.710 42.015 10.730 ;
        RECT 46.365 10.710 47.015 10.730 ;
        RECT 51.365 10.710 52.015 10.730 ;
        RECT 4.785 10.440 7.015 10.710 ;
        RECT 9.785 10.440 12.015 10.710 ;
        RECT 14.785 10.440 17.015 10.710 ;
        RECT 19.785 10.440 22.015 10.710 ;
        RECT 24.785 10.440 27.015 10.710 ;
        RECT 29.785 10.440 32.015 10.710 ;
        RECT 34.785 10.440 37.015 10.710 ;
        RECT 39.785 10.440 42.015 10.710 ;
        RECT 44.785 10.440 47.015 10.710 ;
        RECT 49.785 10.440 52.015 10.710 ;
        RECT 4.785 10.375 7.005 10.440 ;
        RECT 9.785 10.375 12.005 10.440 ;
        RECT 14.785 10.375 17.005 10.440 ;
        RECT 19.785 10.375 22.005 10.440 ;
        RECT 24.785 10.375 27.005 10.440 ;
        RECT 29.785 10.375 32.005 10.440 ;
        RECT 34.785 10.375 37.005 10.440 ;
        RECT 39.785 10.375 42.005 10.440 ;
        RECT 44.785 10.375 47.005 10.440 ;
        RECT 49.785 10.375 52.005 10.440 ;
        RECT 4.785 9.580 5.410 10.375 ;
        RECT 9.785 9.580 10.410 10.375 ;
        RECT 14.785 9.580 15.410 10.375 ;
        RECT 19.785 9.580 20.410 10.375 ;
        RECT 24.785 9.580 25.410 10.375 ;
        RECT 29.785 9.580 30.410 10.375 ;
        RECT 34.785 9.580 35.410 10.375 ;
        RECT 39.785 9.580 40.410 10.375 ;
        RECT 44.785 9.580 45.410 10.375 ;
        RECT 49.785 9.580 50.410 10.375 ;
        RECT 4.785 8.580 5.640 9.580 ;
        RECT 9.785 8.580 10.640 9.580 ;
        RECT 14.785 8.580 15.640 9.580 ;
        RECT 19.785 8.580 20.640 9.580 ;
        RECT 24.785 8.580 25.640 9.580 ;
        RECT 29.785 8.580 30.640 9.580 ;
        RECT 34.785 8.580 35.640 9.580 ;
        RECT 39.785 8.580 40.640 9.580 ;
        RECT 44.785 8.580 45.640 9.580 ;
        RECT 49.785 8.580 50.640 9.580 ;
        RECT 4.785 7.080 5.410 8.580 ;
        RECT 9.785 7.080 10.410 8.580 ;
        RECT 14.785 7.080 15.410 8.580 ;
        RECT 19.785 7.080 20.410 8.580 ;
        RECT 24.785 7.080 25.410 8.580 ;
        RECT 29.785 7.080 30.410 8.580 ;
        RECT 34.785 7.080 35.410 8.580 ;
        RECT 39.785 7.080 40.410 8.580 ;
        RECT 44.785 7.080 45.410 8.580 ;
        RECT 49.785 7.080 50.410 8.580 ;
        RECT 4.785 6.080 5.640 7.080 ;
        RECT 9.785 6.080 10.640 7.080 ;
        RECT 14.785 6.080 15.640 7.080 ;
        RECT 19.785 6.080 20.640 7.080 ;
        RECT 24.785 6.080 25.640 7.080 ;
        RECT 29.785 6.080 30.640 7.080 ;
        RECT 34.785 6.080 35.640 7.080 ;
        RECT 39.785 6.080 40.640 7.080 ;
        RECT 44.785 6.080 45.640 7.080 ;
        RECT 49.785 6.080 50.640 7.080 ;
        RECT 4.785 5.050 5.410 6.080 ;
        RECT 9.785 5.050 10.410 6.080 ;
        RECT 14.785 5.050 15.410 6.080 ;
        RECT 19.785 5.050 20.410 6.080 ;
        RECT 24.785 5.050 25.410 6.080 ;
        RECT 29.785 5.050 30.410 6.080 ;
        RECT 34.785 5.050 35.410 6.080 ;
        RECT 39.785 5.050 40.410 6.080 ;
        RECT 44.785 5.050 45.410 6.080 ;
        RECT 49.785 5.050 50.410 6.080 ;
        RECT 4.785 5.045 7.005 5.050 ;
        RECT 9.785 5.045 12.005 5.050 ;
        RECT 14.785 5.045 17.005 5.050 ;
        RECT 19.785 5.045 22.005 5.050 ;
        RECT 24.785 5.045 27.005 5.050 ;
        RECT 29.785 5.045 32.005 5.050 ;
        RECT 34.785 5.045 37.005 5.050 ;
        RECT 39.785 5.045 42.005 5.050 ;
        RECT 44.785 5.045 47.005 5.050 ;
        RECT 49.785 5.045 52.005 5.050 ;
        RECT 4.785 4.755 7.010 5.045 ;
        RECT 9.785 4.755 12.010 5.045 ;
        RECT 14.785 4.755 17.010 5.045 ;
        RECT 19.785 4.755 22.010 5.045 ;
        RECT 24.785 4.755 27.010 5.045 ;
        RECT 29.785 4.755 32.010 5.045 ;
        RECT 34.785 4.755 37.010 5.045 ;
        RECT 39.785 4.755 42.010 5.045 ;
        RECT 44.785 4.755 47.010 5.045 ;
        RECT 49.785 4.755 52.010 5.045 ;
        RECT 4.785 4.715 7.005 4.755 ;
        RECT 9.785 4.715 12.005 4.755 ;
        RECT 14.785 4.715 17.005 4.755 ;
        RECT 19.785 4.715 22.005 4.755 ;
        RECT 24.785 4.715 27.005 4.755 ;
        RECT 29.785 4.715 32.005 4.755 ;
        RECT 34.785 4.715 37.005 4.755 ;
        RECT 39.785 4.715 42.005 4.755 ;
        RECT 44.785 4.715 47.005 4.755 ;
        RECT 49.785 4.715 52.005 4.755 ;
        RECT 4.785 3.565 5.410 4.715 ;
        RECT 9.785 3.565 10.410 4.715 ;
        RECT 14.785 3.565 15.410 4.715 ;
        RECT 19.785 3.565 20.410 4.715 ;
        RECT 24.785 3.565 25.410 4.715 ;
        RECT 29.785 3.565 30.410 4.715 ;
        RECT 34.785 3.565 35.410 4.715 ;
        RECT 39.785 3.565 40.410 4.715 ;
        RECT 44.785 3.565 45.410 4.715 ;
        RECT 49.785 3.565 50.410 4.715 ;
        RECT -45.995 2.475 54.090 3.565 ;
      LAYER via ;
        RECT -23.840 29.450 -23.580 29.710 ;
        RECT -23.840 29.130 -23.580 29.390 ;
        RECT 105.445 29.650 105.705 29.910 ;
        RECT 105.445 29.330 105.705 29.590 ;
        RECT -23.835 13.495 -23.575 13.755 ;
        RECT -23.835 13.175 -23.575 13.435 ;
        RECT -23.835 3.060 -23.575 3.320 ;
        RECT -23.835 2.740 -23.575 3.000 ;
      LAYER met2 ;
        RECT 105.415 29.765 105.735 29.940 ;
        RECT -23.970 29.265 105.775 29.765 ;
        RECT -23.870 29.100 -23.550 29.265 ;
        RECT -23.900 2.535 -23.510 13.810 ;
    END
  END vss
  PIN bias
    ANTENNAGATEAREA 40.000000 ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER li1 ;
        RECT 5.670 9.770 7.670 9.940 ;
        RECT 10.670 9.770 12.670 9.940 ;
        RECT 15.670 9.770 17.670 9.940 ;
        RECT 20.670 9.770 22.670 9.940 ;
        RECT 25.670 9.770 27.670 9.940 ;
        RECT 30.670 9.770 32.670 9.940 ;
        RECT 35.670 9.770 37.670 9.940 ;
        RECT 40.670 9.770 42.670 9.940 ;
        RECT 45.670 9.770 47.670 9.940 ;
        RECT 50.670 9.770 52.670 9.940 ;
        RECT 7.730 8.560 7.900 9.600 ;
        RECT 5.670 8.220 7.670 8.390 ;
        RECT 10.670 8.220 12.670 8.390 ;
        RECT 15.670 8.220 17.670 8.390 ;
        RECT 20.670 8.220 22.670 8.390 ;
        RECT 25.670 8.220 27.670 8.390 ;
        RECT 30.670 8.220 32.670 8.390 ;
        RECT 35.670 8.220 37.670 8.390 ;
        RECT 40.670 8.220 42.670 8.390 ;
        RECT 45.670 8.220 47.670 8.390 ;
        RECT 50.670 8.220 52.670 8.390 ;
        RECT 5.670 7.270 7.670 7.440 ;
        RECT 10.670 7.270 12.670 7.440 ;
        RECT 15.670 7.270 17.670 7.440 ;
        RECT 20.670 7.270 22.670 7.440 ;
        RECT 25.670 7.270 27.670 7.440 ;
        RECT 30.670 7.270 32.670 7.440 ;
        RECT 35.670 7.270 37.670 7.440 ;
        RECT 40.670 7.270 42.670 7.440 ;
        RECT 45.670 7.270 47.670 7.440 ;
        RECT 50.670 7.270 52.670 7.440 ;
        RECT 7.730 6.060 7.900 7.100 ;
        RECT 5.670 5.720 7.670 5.890 ;
        RECT 10.670 5.720 12.670 5.890 ;
        RECT 15.670 5.720 17.670 5.890 ;
        RECT 20.670 5.720 22.670 5.890 ;
        RECT 25.670 5.720 27.670 5.890 ;
        RECT 30.670 5.720 32.670 5.890 ;
        RECT 35.670 5.720 37.670 5.890 ;
        RECT 40.670 5.720 42.670 5.890 ;
        RECT 45.670 5.720 47.670 5.890 ;
        RECT 50.670 5.720 52.670 5.890 ;
      LAYER met1 ;
        RECT -45.995 11.435 8.555 12.055 ;
        RECT 5.690 9.740 7.650 9.970 ;
        RECT 7.930 9.580 8.555 11.435 ;
        RECT 10.690 9.740 12.650 9.970 ;
        RECT 15.690 9.740 17.650 9.970 ;
        RECT 20.690 9.740 22.650 9.970 ;
        RECT 25.690 9.740 27.650 9.970 ;
        RECT 30.690 9.740 32.650 9.970 ;
        RECT 35.690 9.740 37.650 9.970 ;
        RECT 40.690 9.740 42.650 9.970 ;
        RECT 45.690 9.740 47.650 9.970 ;
        RECT 50.690 9.740 52.650 9.970 ;
        RECT 7.700 8.580 8.555 9.580 ;
        RECT 5.690 8.185 7.650 8.420 ;
        RECT 7.930 8.185 8.555 8.580 ;
        RECT 5.690 7.465 8.555 8.185 ;
        RECT 5.690 7.240 7.650 7.465 ;
        RECT 7.930 7.080 8.555 7.465 ;
        RECT 10.690 7.240 12.650 8.420 ;
        RECT 15.690 7.240 17.650 8.420 ;
        RECT 20.690 7.240 22.650 8.420 ;
        RECT 25.690 7.240 27.650 8.420 ;
        RECT 30.690 7.240 32.650 8.420 ;
        RECT 35.690 7.240 37.650 8.420 ;
        RECT 40.690 7.240 42.650 8.420 ;
        RECT 45.690 7.240 47.650 8.420 ;
        RECT 50.690 7.240 52.650 8.420 ;
        RECT 7.700 6.080 8.555 7.080 ;
        RECT 5.690 5.690 7.650 5.920 ;
        RECT 7.930 4.300 8.555 6.080 ;
        RECT 10.690 5.690 12.650 5.920 ;
        RECT 15.690 5.690 17.650 5.920 ;
        RECT 20.690 5.690 22.650 5.920 ;
        RECT 25.690 5.690 27.650 5.920 ;
        RECT 30.690 5.690 32.650 5.920 ;
        RECT 35.690 5.690 37.650 5.920 ;
        RECT 40.690 5.690 42.650 5.920 ;
        RECT 45.690 5.690 47.650 5.920 ;
        RECT 50.690 5.690 52.650 5.920 ;
      LAYER via ;
        RECT 6.415 7.705 6.675 7.965 ;
        RECT 6.735 7.705 6.995 7.965 ;
        RECT 11.415 7.705 11.675 7.965 ;
        RECT 11.735 7.705 11.995 7.965 ;
        RECT 16.415 7.705 16.675 7.965 ;
        RECT 16.735 7.705 16.995 7.965 ;
        RECT 21.415 7.705 21.675 7.965 ;
        RECT 21.735 7.705 21.995 7.965 ;
        RECT 26.415 7.705 26.675 7.965 ;
        RECT 26.735 7.705 26.995 7.965 ;
        RECT 31.415 7.705 31.675 7.965 ;
        RECT 31.735 7.705 31.995 7.965 ;
        RECT 36.415 7.705 36.675 7.965 ;
        RECT 36.735 7.705 36.995 7.965 ;
        RECT 41.415 7.705 41.675 7.965 ;
        RECT 41.735 7.705 41.995 7.965 ;
        RECT 46.415 7.705 46.675 7.965 ;
        RECT 46.735 7.705 46.995 7.965 ;
        RECT 51.415 7.705 51.675 7.965 ;
        RECT 51.735 7.705 51.995 7.965 ;
      LAYER met2 ;
        RECT 6.340 7.625 52.135 8.045 ;
    END
  END bias
  PIN vdd
    ANTENNADIFFAREA 11.599999 ;
    PORT
      LAYER li1 ;
        RECT 10.755 43.520 11.445 43.850 ;
        RECT 15.755 43.520 16.445 43.850 ;
        RECT 9.890 40.525 10.060 42.565 ;
        RECT 14.890 40.525 15.060 42.565 ;
        RECT 9.890 36.825 10.060 38.865 ;
        RECT 14.890 36.825 15.060 38.865 ;
        RECT 10.740 35.495 11.430 35.825 ;
        RECT 15.740 35.495 16.430 35.825 ;
        RECT 59.345 35.220 60.035 35.550 ;
        RECT 63.845 35.220 64.535 35.550 ;
        RECT 68.345 35.220 69.035 35.550 ;
        RECT 72.845 35.220 73.535 35.550 ;
        RECT 77.345 35.220 78.035 35.550 ;
        RECT 81.845 35.220 82.535 35.550 ;
        RECT 86.345 35.220 87.035 35.550 ;
        RECT 90.845 35.220 91.535 35.550 ;
        RECT 58.480 32.225 58.650 34.265 ;
        RECT 62.980 32.225 63.150 34.265 ;
        RECT 67.480 32.225 67.650 34.265 ;
        RECT 71.980 32.225 72.150 34.265 ;
        RECT 76.480 32.225 76.650 34.265 ;
        RECT 80.980 32.225 81.150 34.265 ;
        RECT 85.480 32.225 85.650 34.265 ;
        RECT 89.980 32.225 90.150 34.265 ;
        RECT 58.480 28.525 58.650 30.565 ;
        RECT 62.980 28.525 63.150 30.565 ;
        RECT 67.480 28.525 67.650 30.565 ;
        RECT 71.980 28.525 72.150 30.565 ;
        RECT 76.480 28.525 76.650 30.565 ;
        RECT 80.980 28.525 81.150 30.565 ;
        RECT 85.480 28.525 85.650 30.565 ;
        RECT 89.980 28.525 90.150 30.565 ;
        RECT 59.330 27.195 60.020 27.525 ;
        RECT 63.830 27.195 64.520 27.525 ;
        RECT 68.330 27.195 69.020 27.525 ;
        RECT 72.830 27.195 73.520 27.525 ;
        RECT 77.330 27.195 78.020 27.525 ;
        RECT 81.830 27.195 82.520 27.525 ;
        RECT 86.330 27.195 87.020 27.525 ;
        RECT 90.830 27.195 91.520 27.525 ;
      LAYER met1 ;
        RECT -45.995 44.755 21.330 45.350 ;
        RECT 9.195 43.945 9.860 44.755 ;
        RECT 14.195 43.945 14.860 44.755 ;
        RECT 9.195 43.425 11.500 43.945 ;
        RECT 14.195 43.425 16.500 43.945 ;
        RECT 9.195 42.545 9.860 43.425 ;
        RECT 14.195 42.545 14.860 43.425 ;
        RECT 9.195 40.545 10.090 42.545 ;
        RECT 14.195 40.545 15.090 42.545 ;
        RECT 9.195 38.845 9.860 40.545 ;
        RECT 14.195 38.845 14.860 40.545 ;
        RECT 9.195 36.845 10.090 38.845 ;
        RECT 14.195 36.845 15.090 38.845 ;
        RECT 20.625 37.370 21.330 44.755 ;
        RECT 9.195 35.920 9.860 36.845 ;
        RECT 14.195 35.920 14.860 36.845 ;
        RECT 20.625 36.455 89.950 37.370 ;
        RECT 9.195 35.400 11.500 35.920 ;
        RECT 14.195 35.400 16.500 35.920 ;
        RECT 57.785 35.645 58.450 36.455 ;
        RECT 62.285 35.645 62.950 36.455 ;
        RECT 66.785 35.645 67.450 36.455 ;
        RECT 71.285 35.645 71.950 36.455 ;
        RECT 75.785 35.645 76.450 36.455 ;
        RECT 80.285 35.645 80.950 36.455 ;
        RECT 84.785 35.645 85.450 36.455 ;
        RECT 89.285 35.645 89.950 36.455 ;
        RECT 57.785 35.125 60.090 35.645 ;
        RECT 62.285 35.125 64.590 35.645 ;
        RECT 66.785 35.125 69.090 35.645 ;
        RECT 71.285 35.125 73.590 35.645 ;
        RECT 75.785 35.125 78.090 35.645 ;
        RECT 80.285 35.125 82.590 35.645 ;
        RECT 84.785 35.125 87.090 35.645 ;
        RECT 89.285 35.125 91.590 35.645 ;
        RECT 57.785 34.245 58.450 35.125 ;
        RECT 62.285 34.245 62.950 35.125 ;
        RECT 66.785 34.245 67.450 35.125 ;
        RECT 71.285 34.245 71.950 35.125 ;
        RECT 75.785 34.245 76.450 35.125 ;
        RECT 80.285 34.245 80.950 35.125 ;
        RECT 84.785 34.245 85.450 35.125 ;
        RECT 89.285 34.245 89.950 35.125 ;
        RECT 57.785 32.245 58.680 34.245 ;
        RECT 62.285 32.245 63.180 34.245 ;
        RECT 66.785 32.245 67.680 34.245 ;
        RECT 71.285 32.245 72.180 34.245 ;
        RECT 75.785 32.245 76.680 34.245 ;
        RECT 80.285 32.245 81.180 34.245 ;
        RECT 84.785 32.245 85.680 34.245 ;
        RECT 89.285 32.245 90.180 34.245 ;
        RECT 57.785 30.545 58.450 32.245 ;
        RECT 62.285 30.545 62.950 32.245 ;
        RECT 66.785 30.545 67.450 32.245 ;
        RECT 71.285 30.545 71.950 32.245 ;
        RECT 75.785 30.545 76.450 32.245 ;
        RECT 80.285 30.545 80.950 32.245 ;
        RECT 84.785 30.545 85.450 32.245 ;
        RECT 89.285 30.545 89.950 32.245 ;
        RECT 57.785 28.545 58.680 30.545 ;
        RECT 62.285 28.545 63.180 30.545 ;
        RECT 66.785 28.545 67.680 30.545 ;
        RECT 71.285 28.545 72.180 30.545 ;
        RECT 75.785 28.545 76.680 30.545 ;
        RECT 80.285 28.545 81.180 30.545 ;
        RECT 84.785 28.545 85.680 30.545 ;
        RECT 89.285 28.545 90.180 30.545 ;
        RECT 57.785 27.620 58.450 28.545 ;
        RECT 62.285 27.620 62.950 28.545 ;
        RECT 66.785 27.620 67.450 28.545 ;
        RECT 71.285 27.620 71.950 28.545 ;
        RECT 75.785 27.620 76.450 28.545 ;
        RECT 80.285 27.620 80.950 28.545 ;
        RECT 84.785 27.620 85.450 28.545 ;
        RECT 89.285 27.620 89.950 28.545 ;
        RECT 57.785 27.100 60.090 27.620 ;
        RECT 62.285 27.100 64.590 27.620 ;
        RECT 66.785 27.100 69.090 27.620 ;
        RECT 71.285 27.100 73.590 27.620 ;
        RECT 75.785 27.100 78.090 27.620 ;
        RECT 80.285 27.100 82.590 27.620 ;
        RECT 84.785 27.100 87.090 27.620 ;
        RECT 89.285 27.100 91.590 27.620 ;
    END
  END vdd
  PIN out
    ANTENNADIFFAREA 13.920000 ;
    PORT
      LAYER li1 ;
        RECT 60.770 32.225 60.940 34.265 ;
        RECT 65.270 32.225 65.440 34.265 ;
        RECT 69.770 32.225 69.940 34.265 ;
        RECT 74.270 32.225 74.440 34.265 ;
        RECT 78.770 32.225 78.940 34.265 ;
        RECT 83.270 32.225 83.440 34.265 ;
        RECT 87.770 32.225 87.940 34.265 ;
        RECT 92.270 32.225 92.440 34.265 ;
        RECT 60.770 28.525 60.940 30.565 ;
        RECT 65.270 28.525 65.440 30.565 ;
        RECT 69.770 28.525 69.940 30.565 ;
        RECT 74.270 28.525 74.440 30.565 ;
        RECT 78.770 28.525 78.940 30.565 ;
        RECT 83.270 28.525 83.440 30.565 ;
        RECT 87.770 28.525 87.940 30.565 ;
        RECT 92.270 28.525 92.440 30.565 ;
        RECT 107.195 30.280 107.885 32.440 ;
        RECT 17.730 8.560 17.900 9.600 ;
        RECT 22.730 8.560 22.900 9.600 ;
        RECT 27.730 8.560 27.900 9.600 ;
        RECT 32.730 8.560 32.900 9.600 ;
        RECT 37.730 8.560 37.900 9.600 ;
        RECT 42.730 8.560 42.900 9.600 ;
        RECT 47.730 8.560 47.900 9.600 ;
        RECT 52.730 8.560 52.900 9.600 ;
        RECT 17.730 6.060 17.900 7.100 ;
        RECT 22.730 6.060 22.900 7.100 ;
        RECT 27.730 6.060 27.900 7.100 ;
        RECT 32.730 6.060 32.900 7.100 ;
        RECT 37.730 6.060 37.900 7.100 ;
        RECT 42.730 6.060 42.900 7.100 ;
        RECT 47.730 6.060 47.900 7.100 ;
        RECT 52.730 6.060 52.900 7.100 ;
      LAYER met1 ;
        RECT 60.970 34.245 61.635 34.900 ;
        RECT 65.470 34.245 66.135 34.900 ;
        RECT 69.970 34.245 70.635 34.900 ;
        RECT 74.470 34.245 75.135 34.900 ;
        RECT 78.970 34.245 79.635 34.900 ;
        RECT 83.470 34.245 84.135 34.900 ;
        RECT 87.970 34.245 88.635 34.900 ;
        RECT 92.470 34.245 93.135 34.900 ;
        RECT 60.740 32.245 61.635 34.245 ;
        RECT 65.240 32.245 66.135 34.245 ;
        RECT 69.740 32.245 70.635 34.245 ;
        RECT 74.240 32.245 75.135 34.245 ;
        RECT 78.740 32.245 79.635 34.245 ;
        RECT 83.240 32.245 84.135 34.245 ;
        RECT 87.740 32.245 88.635 34.245 ;
        RECT 92.240 32.245 93.135 34.245 ;
        RECT 60.970 30.545 61.635 32.245 ;
        RECT 65.470 30.545 66.135 32.245 ;
        RECT 69.970 30.545 70.635 32.245 ;
        RECT 74.470 30.545 75.135 32.245 ;
        RECT 78.970 30.545 79.635 32.245 ;
        RECT 83.470 30.545 84.135 32.245 ;
        RECT 87.970 30.545 88.635 32.245 ;
        RECT 92.470 30.545 93.135 32.245 ;
        RECT 60.740 28.545 61.635 30.545 ;
        RECT 65.240 28.545 66.135 30.545 ;
        RECT 69.740 28.545 70.635 30.545 ;
        RECT 74.240 28.545 75.135 30.545 ;
        RECT 78.740 28.545 79.635 30.545 ;
        RECT 83.240 28.545 84.135 30.545 ;
        RECT 87.740 28.545 88.635 30.545 ;
        RECT 92.240 28.545 93.135 30.545 ;
        RECT 60.970 26.250 61.635 28.545 ;
        RECT 65.470 26.250 66.135 28.545 ;
        RECT 69.970 26.250 70.635 28.545 ;
        RECT 74.470 26.250 75.135 28.545 ;
        RECT 78.970 26.250 79.635 28.545 ;
        RECT 83.470 26.250 84.135 28.545 ;
        RECT 87.970 26.250 88.635 28.545 ;
        RECT 92.470 26.250 93.135 28.545 ;
        RECT 60.970 25.320 93.135 26.250 ;
        RECT 61.455 19.875 62.305 25.320 ;
        RECT 107.245 19.875 107.835 32.415 ;
        RECT 61.455 18.695 169.250 19.875 ;
        RECT 61.455 12.600 62.305 18.695 ;
        RECT 17.930 11.985 62.305 12.600 ;
        RECT 17.930 9.580 18.555 11.985 ;
        RECT 22.930 9.580 23.555 11.985 ;
        RECT 27.930 9.580 28.555 11.985 ;
        RECT 32.930 9.580 33.555 11.985 ;
        RECT 37.930 9.580 38.555 11.985 ;
        RECT 42.930 9.580 43.555 11.985 ;
        RECT 47.930 9.580 48.555 11.985 ;
        RECT 52.930 9.580 53.555 11.985 ;
        RECT 17.700 8.580 18.555 9.580 ;
        RECT 22.700 8.580 23.555 9.580 ;
        RECT 27.700 8.580 28.555 9.580 ;
        RECT 32.700 8.580 33.555 9.580 ;
        RECT 37.700 8.580 38.555 9.580 ;
        RECT 42.700 8.580 43.555 9.580 ;
        RECT 47.700 8.580 48.555 9.580 ;
        RECT 52.700 8.580 53.555 9.580 ;
        RECT 17.930 7.080 18.555 8.580 ;
        RECT 22.930 7.080 23.555 8.580 ;
        RECT 27.930 7.080 28.555 8.580 ;
        RECT 32.930 7.080 33.555 8.580 ;
        RECT 37.930 7.080 38.555 8.580 ;
        RECT 42.930 7.080 43.555 8.580 ;
        RECT 47.930 7.080 48.555 8.580 ;
        RECT 52.930 7.080 53.555 8.580 ;
        RECT 17.700 6.080 18.555 7.080 ;
        RECT 22.700 6.080 23.555 7.080 ;
        RECT 27.700 6.080 28.555 7.080 ;
        RECT 32.700 6.080 33.555 7.080 ;
        RECT 37.700 6.080 38.555 7.080 ;
        RECT 42.700 6.080 43.555 7.080 ;
        RECT 47.700 6.080 48.555 7.080 ;
        RECT 52.700 6.080 53.555 7.080 ;
        RECT 17.930 4.300 18.555 6.080 ;
        RECT 22.930 4.300 23.555 6.080 ;
        RECT 27.930 4.300 28.555 6.080 ;
        RECT 32.930 4.300 33.555 6.080 ;
        RECT 37.930 4.300 38.555 6.080 ;
        RECT 42.930 4.300 43.555 6.080 ;
        RECT 47.930 4.300 48.555 6.080 ;
        RECT 52.930 4.300 53.555 6.080 ;
    END
  END out
  PIN in_n
    ANTENNAGATEAREA 100.000000 ;
    PORT
      LAYER li1 ;
        RECT -21.040 28.340 -20.040 28.510 ;
        RECT -17.540 28.340 -16.540 28.510 ;
        RECT -14.040 28.340 -13.040 28.510 ;
        RECT -10.540 28.340 -9.540 28.510 ;
        RECT -7.040 28.340 -6.040 28.510 ;
        RECT -3.540 28.340 -2.540 28.510 ;
        RECT -0.040 28.340 0.960 28.510 ;
        RECT 3.460 28.340 4.460 28.510 ;
        RECT 6.960 28.340 7.960 28.510 ;
        RECT 10.460 28.340 11.460 28.510 ;
        RECT -21.040 17.790 -20.040 17.960 ;
        RECT -17.540 17.790 -16.540 17.960 ;
        RECT -14.040 17.790 -13.040 17.960 ;
        RECT -10.540 17.790 -9.540 17.960 ;
        RECT -7.040 17.790 -6.040 17.960 ;
        RECT -3.540 17.790 -2.540 17.960 ;
        RECT -0.040 17.790 0.960 17.960 ;
        RECT 3.460 17.790 4.460 17.960 ;
        RECT 6.960 17.790 7.960 17.960 ;
        RECT 10.460 17.790 11.460 17.960 ;
      LAYER met1 ;
        RECT -21.020 28.310 -20.060 28.540 ;
        RECT -17.520 28.310 -16.560 28.540 ;
        RECT -14.020 28.310 -13.060 28.540 ;
        RECT -10.520 28.310 -9.560 28.540 ;
        RECT -7.020 28.310 -6.060 28.540 ;
        RECT -3.520 28.310 -2.560 28.540 ;
        RECT -0.020 28.310 0.940 28.540 ;
        RECT 3.480 28.310 4.440 28.540 ;
        RECT 6.980 28.310 7.940 28.540 ;
        RECT 10.480 28.310 11.440 28.540 ;
        RECT -21.020 16.785 -20.060 17.990 ;
        RECT -17.520 16.785 -16.560 17.990 ;
        RECT -14.020 16.785 -13.060 17.990 ;
        RECT -10.520 16.785 -9.560 17.990 ;
        RECT -7.020 16.785 -6.060 17.990 ;
        RECT -3.520 16.785 -2.560 17.990 ;
        RECT -0.020 16.785 0.940 17.990 ;
        RECT 3.480 16.785 4.440 17.990 ;
        RECT 6.980 16.785 7.940 17.990 ;
        RECT 10.480 16.785 11.440 17.990 ;
      LAYER via ;
        RECT -20.825 17.155 -20.565 17.415 ;
        RECT -20.505 17.155 -20.245 17.415 ;
        RECT -17.325 17.155 -17.065 17.415 ;
        RECT -17.005 17.155 -16.745 17.415 ;
        RECT -13.825 17.155 -13.565 17.415 ;
        RECT -13.505 17.155 -13.245 17.415 ;
        RECT -10.325 17.155 -10.065 17.415 ;
        RECT -10.005 17.155 -9.745 17.415 ;
        RECT -6.825 17.155 -6.565 17.415 ;
        RECT -6.505 17.155 -6.245 17.415 ;
        RECT -3.325 17.155 -3.065 17.415 ;
        RECT -3.005 17.155 -2.745 17.415 ;
        RECT 0.175 17.155 0.435 17.415 ;
        RECT 0.495 17.155 0.755 17.415 ;
        RECT 3.675 17.155 3.935 17.415 ;
        RECT 3.995 17.155 4.255 17.415 ;
        RECT 7.175 17.155 7.435 17.415 ;
        RECT 7.495 17.155 7.755 17.415 ;
        RECT 10.675 17.155 10.935 17.415 ;
        RECT 10.995 17.155 11.255 17.415 ;
      LAYER met2 ;
        RECT -45.995 17.070 11.365 17.495 ;
    END
  END in_n
  PIN in_p
    ANTENNAGATEAREA 100.000000 ;
    PORT
      LAYER li1 ;
        RECT 18.960 28.340 19.960 28.510 ;
        RECT 22.460 28.340 23.460 28.510 ;
        RECT 25.960 28.340 26.960 28.510 ;
        RECT 29.460 28.340 30.460 28.510 ;
        RECT 32.960 28.340 33.960 28.510 ;
        RECT 36.460 28.340 37.460 28.510 ;
        RECT 39.960 28.340 40.960 28.510 ;
        RECT 43.460 28.340 44.460 28.510 ;
        RECT 46.960 28.340 47.960 28.510 ;
        RECT 50.460 28.340 51.460 28.510 ;
        RECT 18.960 17.790 19.960 17.960 ;
        RECT 22.460 17.790 23.460 17.960 ;
        RECT 25.960 17.790 26.960 17.960 ;
        RECT 29.460 17.790 30.460 17.960 ;
        RECT 32.960 17.790 33.960 17.960 ;
        RECT 36.460 17.790 37.460 17.960 ;
        RECT 39.960 17.790 40.960 17.960 ;
        RECT 43.460 17.790 44.460 17.960 ;
        RECT 46.960 17.790 47.960 17.960 ;
        RECT 50.460 17.790 51.460 17.960 ;
      LAYER met1 ;
        RECT 18.980 28.310 19.940 28.540 ;
        RECT 22.480 28.310 23.440 28.540 ;
        RECT 25.980 28.310 26.940 28.540 ;
        RECT 29.480 28.310 30.440 28.540 ;
        RECT 32.980 28.310 33.940 28.540 ;
        RECT 36.480 28.310 37.440 28.540 ;
        RECT 39.980 28.310 40.940 28.540 ;
        RECT 43.480 28.310 44.440 28.540 ;
        RECT 46.980 28.310 47.940 28.540 ;
        RECT 50.480 28.310 51.440 28.540 ;
        RECT 18.980 16.785 19.940 17.990 ;
        RECT 22.480 16.785 23.440 17.990 ;
        RECT 25.980 16.785 26.940 17.990 ;
        RECT 29.480 16.785 30.440 17.990 ;
        RECT 32.980 16.785 33.940 17.990 ;
        RECT 36.480 16.785 37.440 17.990 ;
        RECT 39.980 16.785 40.940 17.990 ;
        RECT 43.480 16.785 44.440 17.990 ;
        RECT 46.980 16.785 47.940 17.990 ;
        RECT 50.480 16.785 51.440 17.990 ;
      LAYER via ;
        RECT 19.175 17.155 19.435 17.415 ;
        RECT 19.495 17.155 19.755 17.415 ;
        RECT 22.675 17.155 22.935 17.415 ;
        RECT 22.995 17.155 23.255 17.415 ;
        RECT 26.175 17.155 26.435 17.415 ;
        RECT 26.495 17.155 26.755 17.415 ;
        RECT 29.675 17.155 29.935 17.415 ;
        RECT 29.995 17.155 30.255 17.415 ;
        RECT 33.175 17.155 33.435 17.415 ;
        RECT 33.495 17.155 33.755 17.415 ;
        RECT 36.675 17.155 36.935 17.415 ;
        RECT 36.995 17.155 37.255 17.415 ;
        RECT 40.175 17.155 40.435 17.415 ;
        RECT 40.495 17.155 40.755 17.415 ;
        RECT 43.675 17.155 43.935 17.415 ;
        RECT 43.995 17.155 44.255 17.415 ;
        RECT 47.175 17.155 47.435 17.415 ;
        RECT 47.495 17.155 47.755 17.415 ;
        RECT 50.675 17.155 50.935 17.415 ;
        RECT 50.995 17.155 51.255 17.415 ;
      LAYER met2 ;
        RECT 19.095 17.070 169.250 17.495 ;
    END
  END in_p
  OBS
      LAYER li1 ;
        RECT 10.120 42.780 12.120 42.950 ;
        RECT 15.120 42.780 17.120 42.950 ;
        RECT 12.180 40.525 12.350 42.565 ;
        RECT 17.180 40.525 17.350 42.565 ;
        RECT 107.195 42.440 107.885 44.600 ;
        RECT 10.120 40.140 12.120 40.310 ;
        RECT 15.120 40.140 17.120 40.310 ;
        RECT 10.120 39.080 12.120 39.250 ;
        RECT 15.120 39.080 17.120 39.250 ;
        RECT 12.180 36.825 12.350 38.865 ;
        RECT 17.180 36.825 17.350 38.865 ;
        RECT 10.120 36.440 12.120 36.610 ;
        RECT 15.120 36.440 17.120 36.610 ;
        RECT 58.710 34.480 60.710 34.650 ;
        RECT 63.210 34.480 65.210 34.650 ;
        RECT 67.710 34.480 69.710 34.650 ;
        RECT 72.210 34.480 74.210 34.650 ;
        RECT 76.710 34.480 78.710 34.650 ;
        RECT 81.210 34.480 83.210 34.650 ;
        RECT 85.710 34.480 87.710 34.650 ;
        RECT 90.210 34.480 92.210 34.650 ;
        RECT 58.710 31.840 60.710 32.010 ;
        RECT 63.210 31.840 65.210 32.010 ;
        RECT 67.710 31.840 69.710 32.010 ;
        RECT 72.210 31.840 74.210 32.010 ;
        RECT 76.710 31.840 78.710 32.010 ;
        RECT 81.210 31.840 83.210 32.010 ;
        RECT 85.710 31.840 87.710 32.010 ;
        RECT 90.210 31.840 92.210 32.010 ;
        RECT 58.710 30.780 60.710 30.950 ;
        RECT 63.210 30.780 65.210 30.950 ;
        RECT 67.710 30.780 69.710 30.950 ;
        RECT 72.210 30.780 74.210 30.950 ;
        RECT 76.710 30.780 78.710 30.950 ;
        RECT 81.210 30.780 83.210 30.950 ;
        RECT 85.710 30.780 87.710 30.950 ;
        RECT 90.210 30.780 92.210 30.950 ;
        RECT -20.840 29.375 -20.150 29.705 ;
        RECT -17.340 29.375 -16.650 29.705 ;
        RECT -13.840 29.375 -13.150 29.705 ;
        RECT -10.340 29.375 -9.650 29.705 ;
        RECT -6.840 29.375 -6.150 29.705 ;
        RECT -3.340 29.375 -2.650 29.705 ;
        RECT 0.160 29.375 0.850 29.705 ;
        RECT 3.660 29.375 4.350 29.705 ;
        RECT 7.160 29.375 7.850 29.705 ;
        RECT 10.660 29.375 11.350 29.705 ;
        RECT 19.160 29.375 19.850 29.705 ;
        RECT 22.660 29.375 23.350 29.705 ;
        RECT 26.160 29.375 26.850 29.705 ;
        RECT 29.660 29.375 30.350 29.705 ;
        RECT 33.160 29.375 33.850 29.705 ;
        RECT 36.660 29.375 37.350 29.705 ;
        RECT 40.160 29.375 40.850 29.705 ;
        RECT 43.660 29.375 44.350 29.705 ;
        RECT 47.160 29.375 47.850 29.705 ;
        RECT 50.660 29.375 51.350 29.705 ;
        RECT -21.270 18.130 -21.100 28.170 ;
        RECT -19.980 18.130 -19.810 28.170 ;
        RECT -17.770 18.130 -17.600 28.170 ;
        RECT -16.480 18.130 -16.310 28.170 ;
        RECT -14.270 18.130 -14.100 28.170 ;
        RECT -12.980 18.130 -12.810 28.170 ;
        RECT -10.770 18.130 -10.600 28.170 ;
        RECT -9.480 18.130 -9.310 28.170 ;
        RECT -7.270 18.130 -7.100 28.170 ;
        RECT -5.980 18.130 -5.810 28.170 ;
        RECT -3.770 18.130 -3.600 28.170 ;
        RECT -2.480 18.130 -2.310 28.170 ;
        RECT -0.270 18.130 -0.100 28.170 ;
        RECT 1.020 18.130 1.190 28.170 ;
        RECT 3.230 18.130 3.400 28.170 ;
        RECT 4.520 18.130 4.690 28.170 ;
        RECT 6.730 18.130 6.900 28.170 ;
        RECT 8.020 18.130 8.190 28.170 ;
        RECT 10.230 18.130 10.400 28.170 ;
        RECT 11.520 18.130 11.690 28.170 ;
        RECT 18.730 18.130 18.900 28.170 ;
        RECT 20.020 18.130 20.190 28.170 ;
        RECT 22.230 18.130 22.400 28.170 ;
        RECT 23.520 18.130 23.690 28.170 ;
        RECT 25.730 18.130 25.900 28.170 ;
        RECT 27.020 18.130 27.190 28.170 ;
        RECT 29.230 18.130 29.400 28.170 ;
        RECT 30.520 18.130 30.690 28.170 ;
        RECT 32.730 18.130 32.900 28.170 ;
        RECT 34.020 18.130 34.190 28.170 ;
        RECT 36.230 18.130 36.400 28.170 ;
        RECT 37.520 18.130 37.690 28.170 ;
        RECT 39.730 18.130 39.900 28.170 ;
        RECT 41.020 18.130 41.190 28.170 ;
        RECT 43.230 18.130 43.400 28.170 ;
        RECT 44.520 18.130 44.690 28.170 ;
        RECT 46.730 18.130 46.900 28.170 ;
        RECT 48.020 18.130 48.190 28.170 ;
        RECT 50.230 18.130 50.400 28.170 ;
        RECT 51.520 18.130 51.690 28.170 ;
        RECT 58.710 28.140 60.710 28.310 ;
        RECT 63.210 28.140 65.210 28.310 ;
        RECT 67.710 28.140 69.710 28.310 ;
        RECT 72.210 28.140 74.210 28.310 ;
        RECT 76.710 28.140 78.710 28.310 ;
        RECT 81.210 28.140 83.210 28.310 ;
        RECT 85.710 28.140 87.710 28.310 ;
        RECT 90.210 28.140 92.210 28.310 ;
        RECT 12.730 8.560 12.900 9.600 ;
        RECT 12.730 6.060 12.900 7.100 ;
      LAYER met1 ;
        RECT 10.140 42.750 12.100 42.980 ;
        RECT 12.380 42.545 13.045 43.200 ;
        RECT 15.140 42.750 17.100 42.980 ;
        RECT 17.380 42.545 18.045 43.200 ;
        RECT 12.150 40.545 13.045 42.545 ;
        RECT 17.150 40.545 18.045 42.545 ;
        RECT 107.245 42.465 107.835 44.570 ;
        RECT 10.140 40.110 12.100 40.340 ;
        RECT 12.380 40.110 13.045 40.545 ;
        RECT 10.140 39.280 13.045 40.110 ;
        RECT 10.140 39.050 12.100 39.280 ;
        RECT 12.380 38.845 13.045 39.280 ;
        RECT 15.140 39.050 17.100 40.340 ;
        RECT 17.380 38.845 18.045 40.545 ;
        RECT 12.150 36.845 13.045 38.845 ;
        RECT 17.150 36.845 18.045 38.845 ;
        RECT 10.140 36.410 12.100 36.640 ;
        RECT 12.380 32.065 13.045 36.845 ;
        RECT 15.140 36.410 17.100 36.640 ;
        RECT 10.060 31.700 13.070 32.065 ;
        RECT 17.380 32.045 18.045 36.845 ;
        RECT 58.730 34.450 60.690 34.680 ;
        RECT 63.230 34.450 65.190 34.680 ;
        RECT 67.730 34.450 69.690 34.680 ;
        RECT 72.230 34.450 74.190 34.680 ;
        RECT 76.730 34.450 78.690 34.680 ;
        RECT 81.230 34.450 83.190 34.680 ;
        RECT 85.730 34.450 87.690 34.680 ;
        RECT 90.230 34.450 92.190 34.680 ;
        RECT -21.980 30.910 13.070 31.700 ;
        RECT 17.385 31.700 18.045 32.045 ;
        RECT 17.385 31.550 50.200 31.700 ;
        RECT 17.385 31.230 50.300 31.550 ;
        RECT 17.385 30.940 50.200 31.230 ;
        RECT -21.980 30.900 10.200 30.910 ;
        RECT -21.980 28.150 -21.300 30.900 ;
        RECT -18.480 28.150 -17.800 30.900 ;
        RECT -14.980 28.150 -14.300 30.900 ;
        RECT -11.480 28.150 -10.800 30.900 ;
        RECT -7.980 28.150 -7.300 30.900 ;
        RECT -4.480 28.150 -3.800 30.900 ;
        RECT -0.980 28.150 -0.300 30.900 ;
        RECT 2.520 28.150 3.200 30.900 ;
        RECT 6.020 28.150 6.700 30.900 ;
        RECT 9.520 28.150 10.200 30.900 ;
        RECT 18.020 30.900 50.200 30.940 ;
        RECT 18.020 28.150 18.700 30.900 ;
        RECT 21.520 28.150 22.200 30.900 ;
        RECT 25.020 28.150 25.700 30.900 ;
        RECT 28.520 28.150 29.200 30.900 ;
        RECT 32.020 28.150 32.700 30.900 ;
        RECT 35.520 28.150 36.200 30.900 ;
        RECT 39.020 28.150 39.700 30.900 ;
        RECT 42.520 28.150 43.200 30.900 ;
        RECT 46.020 28.150 46.700 30.900 ;
        RECT 49.520 28.150 50.200 30.900 ;
        RECT 58.730 30.750 60.690 32.040 ;
        RECT 63.230 30.750 65.190 32.040 ;
        RECT 67.730 30.750 69.690 32.040 ;
        RECT 72.230 30.750 74.190 32.040 ;
        RECT 76.730 30.750 78.690 32.040 ;
        RECT 81.230 30.750 83.190 32.040 ;
        RECT 85.730 30.750 87.690 32.040 ;
        RECT 90.230 30.750 92.190 32.040 ;
        RECT -21.980 18.150 -21.070 28.150 ;
        RECT -20.010 18.150 -19.100 28.150 ;
        RECT -18.480 18.150 -17.570 28.150 ;
        RECT -16.510 18.150 -15.600 28.150 ;
        RECT -14.980 18.150 -14.070 28.150 ;
        RECT -13.010 18.150 -12.100 28.150 ;
        RECT -11.480 18.150 -10.570 28.150 ;
        RECT -9.510 18.150 -8.600 28.150 ;
        RECT -7.980 18.150 -7.070 28.150 ;
        RECT -6.010 18.150 -5.100 28.150 ;
        RECT -4.480 18.150 -3.570 28.150 ;
        RECT -2.510 18.150 -1.600 28.150 ;
        RECT -0.980 18.150 -0.070 28.150 ;
        RECT 0.990 18.150 1.900 28.150 ;
        RECT 2.520 18.150 3.430 28.150 ;
        RECT 4.490 18.150 5.400 28.150 ;
        RECT 6.020 18.150 6.930 28.150 ;
        RECT 7.990 18.150 8.900 28.150 ;
        RECT 9.520 18.150 10.430 28.150 ;
        RECT 11.490 18.150 12.400 28.150 ;
        RECT 18.020 18.150 18.930 28.150 ;
        RECT 19.990 18.150 20.900 28.150 ;
        RECT 21.520 18.150 22.430 28.150 ;
        RECT 23.490 18.150 24.400 28.150 ;
        RECT 25.020 18.150 25.930 28.150 ;
        RECT 26.990 18.150 27.900 28.150 ;
        RECT 28.520 18.150 29.430 28.150 ;
        RECT 30.490 18.150 31.400 28.150 ;
        RECT 32.020 18.150 32.930 28.150 ;
        RECT 33.990 18.150 34.900 28.150 ;
        RECT 35.520 18.150 36.430 28.150 ;
        RECT 37.490 18.150 38.400 28.150 ;
        RECT 39.020 18.150 39.930 28.150 ;
        RECT 40.990 18.150 41.900 28.150 ;
        RECT 42.520 18.150 43.430 28.150 ;
        RECT 44.490 18.150 45.400 28.150 ;
        RECT 46.020 18.150 46.930 28.150 ;
        RECT 47.990 18.150 48.900 28.150 ;
        RECT 49.520 18.150 50.430 28.150 ;
        RECT 51.490 18.150 52.400 28.150 ;
        RECT 58.730 28.110 60.690 28.340 ;
        RECT 63.230 28.110 65.190 28.340 ;
        RECT 67.730 28.110 69.690 28.340 ;
        RECT 72.230 28.110 74.190 28.340 ;
        RECT 76.730 28.110 78.690 28.340 ;
        RECT 81.230 28.110 83.190 28.340 ;
        RECT 85.730 28.110 87.690 28.340 ;
        RECT 90.230 28.110 92.190 28.340 ;
        RECT -19.780 15.400 -19.100 18.150 ;
        RECT -16.280 15.400 -15.600 18.150 ;
        RECT -12.780 15.400 -12.100 18.150 ;
        RECT -9.280 15.400 -8.600 18.150 ;
        RECT -5.780 15.400 -5.100 18.150 ;
        RECT -2.280 15.400 -1.600 18.150 ;
        RECT 1.220 15.400 1.900 18.150 ;
        RECT 4.720 15.400 5.400 18.150 ;
        RECT 8.220 15.400 8.900 18.150 ;
        RECT 11.720 15.400 12.400 18.150 ;
        RECT 20.220 15.400 20.900 18.150 ;
        RECT 23.720 15.400 24.400 18.150 ;
        RECT 27.220 15.400 27.900 18.150 ;
        RECT 30.720 15.400 31.400 18.150 ;
        RECT 34.220 15.400 34.900 18.150 ;
        RECT 37.720 15.400 38.400 18.150 ;
        RECT 41.220 15.400 41.900 18.150 ;
        RECT 44.720 15.400 45.400 18.150 ;
        RECT 48.220 15.400 48.900 18.150 ;
        RECT 51.720 15.400 52.400 18.150 ;
        RECT -19.780 14.600 52.400 15.400 ;
        RECT 12.930 9.580 13.555 14.600 ;
        RECT 12.700 8.580 13.555 9.580 ;
        RECT 12.930 7.080 13.555 8.580 ;
        RECT 12.700 6.080 13.555 7.080 ;
        RECT 12.930 4.300 13.555 6.080 ;
      LAYER via ;
        RECT 107.405 44.175 107.665 44.435 ;
        RECT 107.405 43.855 107.665 44.115 ;
        RECT 10.880 39.585 11.140 39.845 ;
        RECT 11.200 39.585 11.460 39.845 ;
        RECT 15.880 39.585 16.140 39.845 ;
        RECT 16.200 39.585 16.460 39.845 ;
        RECT 49.690 31.260 49.950 31.520 ;
        RECT 50.010 31.260 50.270 31.520 ;
        RECT 59.470 31.265 59.730 31.525 ;
        RECT 59.790 31.265 60.050 31.525 ;
        RECT 63.970 31.265 64.230 31.525 ;
        RECT 64.290 31.265 64.550 31.525 ;
        RECT 68.470 31.265 68.730 31.525 ;
        RECT 68.790 31.265 69.050 31.525 ;
        RECT 72.970 31.265 73.230 31.525 ;
        RECT 73.290 31.265 73.550 31.525 ;
        RECT 77.470 31.265 77.730 31.525 ;
        RECT 77.790 31.265 78.050 31.525 ;
        RECT 81.970 31.265 82.230 31.525 ;
        RECT 82.290 31.265 82.550 31.525 ;
        RECT 86.470 31.265 86.730 31.525 ;
        RECT 86.790 31.265 87.050 31.525 ;
        RECT 90.970 31.265 91.230 31.525 ;
        RECT 91.290 31.265 91.550 31.525 ;
      LAYER met2 ;
        RECT 10.815 39.520 16.515 39.895 ;
        RECT 58.365 31.645 59.190 85.605 ;
        RECT 107.300 43.715 107.780 44.525 ;
        RECT 49.400 31.145 91.655 31.645 ;
      LAYER via2 ;
        RECT 58.630 85.145 58.910 85.425 ;
        RECT 58.630 84.745 58.910 85.025 ;
        RECT 107.390 44.195 107.670 44.475 ;
        RECT 107.390 43.795 107.670 44.075 ;
      LAYER met3 ;
        RECT 58.590 85.535 58.970 85.560 ;
        RECT 58.535 84.625 59.020 85.535 ;
        RECT -43.595 51.845 -12.595 83.340 ;
        RECT -8.595 51.845 22.405 83.340 ;
        RECT 26.405 51.845 57.405 83.340 ;
        RECT 61.405 51.845 92.405 83.340 ;
        RECT 96.405 51.845 127.405 83.340 ;
        RECT 131.405 51.845 162.405 83.340 ;
        RECT 107.350 44.535 107.730 44.580 ;
        RECT 107.290 43.700 107.790 44.535 ;
        RECT 107.350 43.650 107.730 43.700 ;
      LAYER via3 ;
        RECT 58.620 85.210 58.940 85.530 ;
        RECT 58.620 84.660 58.940 84.980 ;
        RECT -43.455 51.945 -43.135 52.265 ;
        RECT -43.055 51.945 -42.735 52.265 ;
        RECT -42.655 51.945 -42.335 52.265 ;
        RECT -42.255 51.945 -41.935 52.265 ;
        RECT -41.855 51.945 -41.535 52.265 ;
        RECT -41.455 51.945 -41.135 52.265 ;
        RECT -41.055 51.945 -40.735 52.265 ;
        RECT -40.655 51.945 -40.335 52.265 ;
        RECT -40.255 51.945 -39.935 52.265 ;
        RECT -39.855 51.945 -39.535 52.265 ;
        RECT -39.455 51.945 -39.135 52.265 ;
        RECT -39.055 51.945 -38.735 52.265 ;
        RECT -38.655 51.945 -38.335 52.265 ;
        RECT -38.255 51.945 -37.935 52.265 ;
        RECT -37.855 51.945 -37.535 52.265 ;
        RECT -37.455 51.945 -37.135 52.265 ;
        RECT -37.055 51.945 -36.735 52.265 ;
        RECT -36.655 51.945 -36.335 52.265 ;
        RECT -36.255 51.945 -35.935 52.265 ;
        RECT -35.855 51.945 -35.535 52.265 ;
        RECT -35.455 51.945 -35.135 52.265 ;
        RECT -35.055 51.945 -34.735 52.265 ;
        RECT -34.655 51.945 -34.335 52.265 ;
        RECT -34.255 51.945 -33.935 52.265 ;
        RECT -33.855 51.945 -33.535 52.265 ;
        RECT -33.455 51.945 -33.135 52.265 ;
        RECT -33.055 51.945 -32.735 52.265 ;
        RECT -32.655 51.945 -32.335 52.265 ;
        RECT -32.255 51.945 -31.935 52.265 ;
        RECT -31.855 51.945 -31.535 52.265 ;
        RECT -31.455 51.945 -31.135 52.265 ;
        RECT -31.055 51.945 -30.735 52.265 ;
        RECT -30.655 51.945 -30.335 52.265 ;
        RECT -30.255 51.945 -29.935 52.265 ;
        RECT -29.855 51.945 -29.535 52.265 ;
        RECT -29.455 51.945 -29.135 52.265 ;
        RECT -29.055 51.945 -28.735 52.265 ;
        RECT -28.655 51.945 -28.335 52.265 ;
        RECT -28.255 51.945 -27.935 52.265 ;
        RECT -27.855 51.945 -27.535 52.265 ;
        RECT -27.455 51.945 -27.135 52.265 ;
        RECT -27.055 51.945 -26.735 52.265 ;
        RECT -26.655 51.945 -26.335 52.265 ;
        RECT -26.255 51.945 -25.935 52.265 ;
        RECT -25.855 51.945 -25.535 52.265 ;
        RECT -25.455 51.945 -25.135 52.265 ;
        RECT -25.055 51.945 -24.735 52.265 ;
        RECT -24.655 51.945 -24.335 52.265 ;
        RECT -24.255 51.945 -23.935 52.265 ;
        RECT -23.855 51.945 -23.535 52.265 ;
        RECT -23.455 51.945 -23.135 52.265 ;
        RECT -23.055 51.945 -22.735 52.265 ;
        RECT -22.655 51.945 -22.335 52.265 ;
        RECT -22.255 51.945 -21.935 52.265 ;
        RECT -21.855 51.945 -21.535 52.265 ;
        RECT -21.455 51.945 -21.135 52.265 ;
        RECT -21.055 51.945 -20.735 52.265 ;
        RECT -20.655 51.945 -20.335 52.265 ;
        RECT -20.255 51.945 -19.935 52.265 ;
        RECT -19.855 51.945 -19.535 52.265 ;
        RECT -19.455 51.945 -19.135 52.265 ;
        RECT -19.055 51.945 -18.735 52.265 ;
        RECT -18.655 51.945 -18.335 52.265 ;
        RECT -18.255 51.945 -17.935 52.265 ;
        RECT -17.855 51.945 -17.535 52.265 ;
        RECT -17.455 51.945 -17.135 52.265 ;
        RECT -17.055 51.945 -16.735 52.265 ;
        RECT -16.655 51.945 -16.335 52.265 ;
        RECT -16.255 51.945 -15.935 52.265 ;
        RECT -15.855 51.945 -15.535 52.265 ;
        RECT -15.455 51.945 -15.135 52.265 ;
        RECT -15.055 51.945 -14.735 52.265 ;
        RECT -14.655 51.945 -14.335 52.265 ;
        RECT -14.255 51.945 -13.935 52.265 ;
        RECT -13.855 51.945 -13.535 52.265 ;
        RECT -13.455 51.945 -13.135 52.265 ;
        RECT -13.055 51.945 -12.735 52.265 ;
        RECT -8.455 51.945 -8.135 52.265 ;
        RECT -8.055 51.945 -7.735 52.265 ;
        RECT -7.655 51.945 -7.335 52.265 ;
        RECT -7.255 51.945 -6.935 52.265 ;
        RECT -6.855 51.945 -6.535 52.265 ;
        RECT -6.455 51.945 -6.135 52.265 ;
        RECT -6.055 51.945 -5.735 52.265 ;
        RECT -5.655 51.945 -5.335 52.265 ;
        RECT -5.255 51.945 -4.935 52.265 ;
        RECT -4.855 51.945 -4.535 52.265 ;
        RECT -4.455 51.945 -4.135 52.265 ;
        RECT -4.055 51.945 -3.735 52.265 ;
        RECT -3.655 51.945 -3.335 52.265 ;
        RECT -3.255 51.945 -2.935 52.265 ;
        RECT -2.855 51.945 -2.535 52.265 ;
        RECT -2.455 51.945 -2.135 52.265 ;
        RECT -2.055 51.945 -1.735 52.265 ;
        RECT -1.655 51.945 -1.335 52.265 ;
        RECT -1.255 51.945 -0.935 52.265 ;
        RECT -0.855 51.945 -0.535 52.265 ;
        RECT -0.455 51.945 -0.135 52.265 ;
        RECT -0.055 51.945 0.265 52.265 ;
        RECT 0.345 51.945 0.665 52.265 ;
        RECT 0.745 51.945 1.065 52.265 ;
        RECT 1.145 51.945 1.465 52.265 ;
        RECT 1.545 51.945 1.865 52.265 ;
        RECT 1.945 51.945 2.265 52.265 ;
        RECT 2.345 51.945 2.665 52.265 ;
        RECT 2.745 51.945 3.065 52.265 ;
        RECT 3.145 51.945 3.465 52.265 ;
        RECT 3.545 51.945 3.865 52.265 ;
        RECT 3.945 51.945 4.265 52.265 ;
        RECT 4.345 51.945 4.665 52.265 ;
        RECT 4.745 51.945 5.065 52.265 ;
        RECT 5.145 51.945 5.465 52.265 ;
        RECT 5.545 51.945 5.865 52.265 ;
        RECT 5.945 51.945 6.265 52.265 ;
        RECT 6.345 51.945 6.665 52.265 ;
        RECT 6.745 51.945 7.065 52.265 ;
        RECT 7.145 51.945 7.465 52.265 ;
        RECT 7.545 51.945 7.865 52.265 ;
        RECT 7.945 51.945 8.265 52.265 ;
        RECT 8.345 51.945 8.665 52.265 ;
        RECT 8.745 51.945 9.065 52.265 ;
        RECT 9.145 51.945 9.465 52.265 ;
        RECT 9.545 51.945 9.865 52.265 ;
        RECT 9.945 51.945 10.265 52.265 ;
        RECT 10.345 51.945 10.665 52.265 ;
        RECT 10.745 51.945 11.065 52.265 ;
        RECT 11.145 51.945 11.465 52.265 ;
        RECT 11.545 51.945 11.865 52.265 ;
        RECT 11.945 51.945 12.265 52.265 ;
        RECT 12.345 51.945 12.665 52.265 ;
        RECT 12.745 51.945 13.065 52.265 ;
        RECT 13.145 51.945 13.465 52.265 ;
        RECT 13.545 51.945 13.865 52.265 ;
        RECT 13.945 51.945 14.265 52.265 ;
        RECT 14.345 51.945 14.665 52.265 ;
        RECT 14.745 51.945 15.065 52.265 ;
        RECT 15.145 51.945 15.465 52.265 ;
        RECT 15.545 51.945 15.865 52.265 ;
        RECT 15.945 51.945 16.265 52.265 ;
        RECT 16.345 51.945 16.665 52.265 ;
        RECT 16.745 51.945 17.065 52.265 ;
        RECT 17.145 51.945 17.465 52.265 ;
        RECT 17.545 51.945 17.865 52.265 ;
        RECT 17.945 51.945 18.265 52.265 ;
        RECT 18.345 51.945 18.665 52.265 ;
        RECT 18.745 51.945 19.065 52.265 ;
        RECT 19.145 51.945 19.465 52.265 ;
        RECT 19.545 51.945 19.865 52.265 ;
        RECT 19.945 51.945 20.265 52.265 ;
        RECT 20.345 51.945 20.665 52.265 ;
        RECT 20.745 51.945 21.065 52.265 ;
        RECT 21.145 51.945 21.465 52.265 ;
        RECT 21.545 51.945 21.865 52.265 ;
        RECT 21.945 51.945 22.265 52.265 ;
        RECT 26.545 51.945 26.865 52.265 ;
        RECT 26.945 51.945 27.265 52.265 ;
        RECT 27.345 51.945 27.665 52.265 ;
        RECT 27.745 51.945 28.065 52.265 ;
        RECT 28.145 51.945 28.465 52.265 ;
        RECT 28.545 51.945 28.865 52.265 ;
        RECT 28.945 51.945 29.265 52.265 ;
        RECT 29.345 51.945 29.665 52.265 ;
        RECT 29.745 51.945 30.065 52.265 ;
        RECT 30.145 51.945 30.465 52.265 ;
        RECT 30.545 51.945 30.865 52.265 ;
        RECT 30.945 51.945 31.265 52.265 ;
        RECT 31.345 51.945 31.665 52.265 ;
        RECT 31.745 51.945 32.065 52.265 ;
        RECT 32.145 51.945 32.465 52.265 ;
        RECT 32.545 51.945 32.865 52.265 ;
        RECT 32.945 51.945 33.265 52.265 ;
        RECT 33.345 51.945 33.665 52.265 ;
        RECT 33.745 51.945 34.065 52.265 ;
        RECT 34.145 51.945 34.465 52.265 ;
        RECT 34.545 51.945 34.865 52.265 ;
        RECT 34.945 51.945 35.265 52.265 ;
        RECT 35.345 51.945 35.665 52.265 ;
        RECT 35.745 51.945 36.065 52.265 ;
        RECT 36.145 51.945 36.465 52.265 ;
        RECT 36.545 51.945 36.865 52.265 ;
        RECT 36.945 51.945 37.265 52.265 ;
        RECT 37.345 51.945 37.665 52.265 ;
        RECT 37.745 51.945 38.065 52.265 ;
        RECT 38.145 51.945 38.465 52.265 ;
        RECT 38.545 51.945 38.865 52.265 ;
        RECT 38.945 51.945 39.265 52.265 ;
        RECT 39.345 51.945 39.665 52.265 ;
        RECT 39.745 51.945 40.065 52.265 ;
        RECT 40.145 51.945 40.465 52.265 ;
        RECT 40.545 51.945 40.865 52.265 ;
        RECT 40.945 51.945 41.265 52.265 ;
        RECT 41.345 51.945 41.665 52.265 ;
        RECT 41.745 51.945 42.065 52.265 ;
        RECT 42.145 51.945 42.465 52.265 ;
        RECT 42.545 51.945 42.865 52.265 ;
        RECT 42.945 51.945 43.265 52.265 ;
        RECT 43.345 51.945 43.665 52.265 ;
        RECT 43.745 51.945 44.065 52.265 ;
        RECT 44.145 51.945 44.465 52.265 ;
        RECT 44.545 51.945 44.865 52.265 ;
        RECT 44.945 51.945 45.265 52.265 ;
        RECT 45.345 51.945 45.665 52.265 ;
        RECT 45.745 51.945 46.065 52.265 ;
        RECT 46.145 51.945 46.465 52.265 ;
        RECT 46.545 51.945 46.865 52.265 ;
        RECT 46.945 51.945 47.265 52.265 ;
        RECT 47.345 51.945 47.665 52.265 ;
        RECT 47.745 51.945 48.065 52.265 ;
        RECT 48.145 51.945 48.465 52.265 ;
        RECT 48.545 51.945 48.865 52.265 ;
        RECT 48.945 51.945 49.265 52.265 ;
        RECT 49.345 51.945 49.665 52.265 ;
        RECT 49.745 51.945 50.065 52.265 ;
        RECT 50.145 51.945 50.465 52.265 ;
        RECT 50.545 51.945 50.865 52.265 ;
        RECT 50.945 51.945 51.265 52.265 ;
        RECT 51.345 51.945 51.665 52.265 ;
        RECT 51.745 51.945 52.065 52.265 ;
        RECT 52.145 51.945 52.465 52.265 ;
        RECT 52.545 51.945 52.865 52.265 ;
        RECT 52.945 51.945 53.265 52.265 ;
        RECT 53.345 51.945 53.665 52.265 ;
        RECT 53.745 51.945 54.065 52.265 ;
        RECT 54.145 51.945 54.465 52.265 ;
        RECT 54.545 51.945 54.865 52.265 ;
        RECT 54.945 51.945 55.265 52.265 ;
        RECT 55.345 51.945 55.665 52.265 ;
        RECT 55.745 51.945 56.065 52.265 ;
        RECT 56.145 51.945 56.465 52.265 ;
        RECT 56.545 51.945 56.865 52.265 ;
        RECT 56.945 51.945 57.265 52.265 ;
        RECT 61.545 51.945 61.865 52.265 ;
        RECT 61.945 51.945 62.265 52.265 ;
        RECT 62.345 51.945 62.665 52.265 ;
        RECT 62.745 51.945 63.065 52.265 ;
        RECT 63.145 51.945 63.465 52.265 ;
        RECT 63.545 51.945 63.865 52.265 ;
        RECT 63.945 51.945 64.265 52.265 ;
        RECT 64.345 51.945 64.665 52.265 ;
        RECT 64.745 51.945 65.065 52.265 ;
        RECT 65.145 51.945 65.465 52.265 ;
        RECT 65.545 51.945 65.865 52.265 ;
        RECT 65.945 51.945 66.265 52.265 ;
        RECT 66.345 51.945 66.665 52.265 ;
        RECT 66.745 51.945 67.065 52.265 ;
        RECT 67.145 51.945 67.465 52.265 ;
        RECT 67.545 51.945 67.865 52.265 ;
        RECT 67.945 51.945 68.265 52.265 ;
        RECT 68.345 51.945 68.665 52.265 ;
        RECT 68.745 51.945 69.065 52.265 ;
        RECT 69.145 51.945 69.465 52.265 ;
        RECT 69.545 51.945 69.865 52.265 ;
        RECT 69.945 51.945 70.265 52.265 ;
        RECT 70.345 51.945 70.665 52.265 ;
        RECT 70.745 51.945 71.065 52.265 ;
        RECT 71.145 51.945 71.465 52.265 ;
        RECT 71.545 51.945 71.865 52.265 ;
        RECT 71.945 51.945 72.265 52.265 ;
        RECT 72.345 51.945 72.665 52.265 ;
        RECT 72.745 51.945 73.065 52.265 ;
        RECT 73.145 51.945 73.465 52.265 ;
        RECT 73.545 51.945 73.865 52.265 ;
        RECT 73.945 51.945 74.265 52.265 ;
        RECT 74.345 51.945 74.665 52.265 ;
        RECT 74.745 51.945 75.065 52.265 ;
        RECT 75.145 51.945 75.465 52.265 ;
        RECT 75.545 51.945 75.865 52.265 ;
        RECT 75.945 51.945 76.265 52.265 ;
        RECT 76.345 51.945 76.665 52.265 ;
        RECT 76.745 51.945 77.065 52.265 ;
        RECT 77.145 51.945 77.465 52.265 ;
        RECT 77.545 51.945 77.865 52.265 ;
        RECT 77.945 51.945 78.265 52.265 ;
        RECT 78.345 51.945 78.665 52.265 ;
        RECT 78.745 51.945 79.065 52.265 ;
        RECT 79.145 51.945 79.465 52.265 ;
        RECT 79.545 51.945 79.865 52.265 ;
        RECT 79.945 51.945 80.265 52.265 ;
        RECT 80.345 51.945 80.665 52.265 ;
        RECT 80.745 51.945 81.065 52.265 ;
        RECT 81.145 51.945 81.465 52.265 ;
        RECT 81.545 51.945 81.865 52.265 ;
        RECT 81.945 51.945 82.265 52.265 ;
        RECT 82.345 51.945 82.665 52.265 ;
        RECT 82.745 51.945 83.065 52.265 ;
        RECT 83.145 51.945 83.465 52.265 ;
        RECT 83.545 51.945 83.865 52.265 ;
        RECT 83.945 51.945 84.265 52.265 ;
        RECT 84.345 51.945 84.665 52.265 ;
        RECT 84.745 51.945 85.065 52.265 ;
        RECT 85.145 51.945 85.465 52.265 ;
        RECT 85.545 51.945 85.865 52.265 ;
        RECT 85.945 51.945 86.265 52.265 ;
        RECT 86.345 51.945 86.665 52.265 ;
        RECT 86.745 51.945 87.065 52.265 ;
        RECT 87.145 51.945 87.465 52.265 ;
        RECT 87.545 51.945 87.865 52.265 ;
        RECT 87.945 51.945 88.265 52.265 ;
        RECT 88.345 51.945 88.665 52.265 ;
        RECT 88.745 51.945 89.065 52.265 ;
        RECT 89.145 51.945 89.465 52.265 ;
        RECT 89.545 51.945 89.865 52.265 ;
        RECT 89.945 51.945 90.265 52.265 ;
        RECT 90.345 51.945 90.665 52.265 ;
        RECT 90.745 51.945 91.065 52.265 ;
        RECT 91.145 51.945 91.465 52.265 ;
        RECT 91.545 51.945 91.865 52.265 ;
        RECT 91.945 51.945 92.265 52.265 ;
        RECT 96.545 51.945 96.865 52.265 ;
        RECT 96.945 51.945 97.265 52.265 ;
        RECT 97.345 51.945 97.665 52.265 ;
        RECT 97.745 51.945 98.065 52.265 ;
        RECT 98.145 51.945 98.465 52.265 ;
        RECT 98.545 51.945 98.865 52.265 ;
        RECT 98.945 51.945 99.265 52.265 ;
        RECT 99.345 51.945 99.665 52.265 ;
        RECT 99.745 51.945 100.065 52.265 ;
        RECT 100.145 51.945 100.465 52.265 ;
        RECT 100.545 51.945 100.865 52.265 ;
        RECT 100.945 51.945 101.265 52.265 ;
        RECT 101.345 51.945 101.665 52.265 ;
        RECT 101.745 51.945 102.065 52.265 ;
        RECT 102.145 51.945 102.465 52.265 ;
        RECT 102.545 51.945 102.865 52.265 ;
        RECT 102.945 51.945 103.265 52.265 ;
        RECT 103.345 51.945 103.665 52.265 ;
        RECT 103.745 51.945 104.065 52.265 ;
        RECT 104.145 51.945 104.465 52.265 ;
        RECT 104.545 51.945 104.865 52.265 ;
        RECT 104.945 51.945 105.265 52.265 ;
        RECT 105.345 51.945 105.665 52.265 ;
        RECT 105.745 51.945 106.065 52.265 ;
        RECT 106.145 51.945 106.465 52.265 ;
        RECT 106.545 51.945 106.865 52.265 ;
        RECT 106.945 51.945 107.265 52.265 ;
        RECT 107.345 51.945 107.665 52.265 ;
        RECT 107.745 51.945 108.065 52.265 ;
        RECT 108.145 51.945 108.465 52.265 ;
        RECT 108.545 51.945 108.865 52.265 ;
        RECT 108.945 51.945 109.265 52.265 ;
        RECT 109.345 51.945 109.665 52.265 ;
        RECT 109.745 51.945 110.065 52.265 ;
        RECT 110.145 51.945 110.465 52.265 ;
        RECT 110.545 51.945 110.865 52.265 ;
        RECT 110.945 51.945 111.265 52.265 ;
        RECT 111.345 51.945 111.665 52.265 ;
        RECT 111.745 51.945 112.065 52.265 ;
        RECT 112.145 51.945 112.465 52.265 ;
        RECT 112.545 51.945 112.865 52.265 ;
        RECT 112.945 51.945 113.265 52.265 ;
        RECT 113.345 51.945 113.665 52.265 ;
        RECT 113.745 51.945 114.065 52.265 ;
        RECT 114.145 51.945 114.465 52.265 ;
        RECT 114.545 51.945 114.865 52.265 ;
        RECT 114.945 51.945 115.265 52.265 ;
        RECT 115.345 51.945 115.665 52.265 ;
        RECT 115.745 51.945 116.065 52.265 ;
        RECT 116.145 51.945 116.465 52.265 ;
        RECT 116.545 51.945 116.865 52.265 ;
        RECT 116.945 51.945 117.265 52.265 ;
        RECT 117.345 51.945 117.665 52.265 ;
        RECT 117.745 51.945 118.065 52.265 ;
        RECT 118.145 51.945 118.465 52.265 ;
        RECT 118.545 51.945 118.865 52.265 ;
        RECT 118.945 51.945 119.265 52.265 ;
        RECT 119.345 51.945 119.665 52.265 ;
        RECT 119.745 51.945 120.065 52.265 ;
        RECT 120.145 51.945 120.465 52.265 ;
        RECT 120.545 51.945 120.865 52.265 ;
        RECT 120.945 51.945 121.265 52.265 ;
        RECT 121.345 51.945 121.665 52.265 ;
        RECT 121.745 51.945 122.065 52.265 ;
        RECT 122.145 51.945 122.465 52.265 ;
        RECT 122.545 51.945 122.865 52.265 ;
        RECT 122.945 51.945 123.265 52.265 ;
        RECT 123.345 51.945 123.665 52.265 ;
        RECT 123.745 51.945 124.065 52.265 ;
        RECT 124.145 51.945 124.465 52.265 ;
        RECT 124.545 51.945 124.865 52.265 ;
        RECT 124.945 51.945 125.265 52.265 ;
        RECT 125.345 51.945 125.665 52.265 ;
        RECT 125.745 51.945 126.065 52.265 ;
        RECT 126.145 51.945 126.465 52.265 ;
        RECT 126.545 51.945 126.865 52.265 ;
        RECT 126.945 51.945 127.265 52.265 ;
        RECT 131.545 51.945 131.865 52.265 ;
        RECT 131.945 51.945 132.265 52.265 ;
        RECT 132.345 51.945 132.665 52.265 ;
        RECT 132.745 51.945 133.065 52.265 ;
        RECT 133.145 51.945 133.465 52.265 ;
        RECT 133.545 51.945 133.865 52.265 ;
        RECT 133.945 51.945 134.265 52.265 ;
        RECT 134.345 51.945 134.665 52.265 ;
        RECT 134.745 51.945 135.065 52.265 ;
        RECT 135.145 51.945 135.465 52.265 ;
        RECT 135.545 51.945 135.865 52.265 ;
        RECT 135.945 51.945 136.265 52.265 ;
        RECT 136.345 51.945 136.665 52.265 ;
        RECT 136.745 51.945 137.065 52.265 ;
        RECT 137.145 51.945 137.465 52.265 ;
        RECT 137.545 51.945 137.865 52.265 ;
        RECT 137.945 51.945 138.265 52.265 ;
        RECT 138.345 51.945 138.665 52.265 ;
        RECT 138.745 51.945 139.065 52.265 ;
        RECT 139.145 51.945 139.465 52.265 ;
        RECT 139.545 51.945 139.865 52.265 ;
        RECT 139.945 51.945 140.265 52.265 ;
        RECT 140.345 51.945 140.665 52.265 ;
        RECT 140.745 51.945 141.065 52.265 ;
        RECT 141.145 51.945 141.465 52.265 ;
        RECT 141.545 51.945 141.865 52.265 ;
        RECT 141.945 51.945 142.265 52.265 ;
        RECT 142.345 51.945 142.665 52.265 ;
        RECT 142.745 51.945 143.065 52.265 ;
        RECT 143.145 51.945 143.465 52.265 ;
        RECT 143.545 51.945 143.865 52.265 ;
        RECT 143.945 51.945 144.265 52.265 ;
        RECT 144.345 51.945 144.665 52.265 ;
        RECT 144.745 51.945 145.065 52.265 ;
        RECT 145.145 51.945 145.465 52.265 ;
        RECT 145.545 51.945 145.865 52.265 ;
        RECT 145.945 51.945 146.265 52.265 ;
        RECT 146.345 51.945 146.665 52.265 ;
        RECT 146.745 51.945 147.065 52.265 ;
        RECT 147.145 51.945 147.465 52.265 ;
        RECT 147.545 51.945 147.865 52.265 ;
        RECT 147.945 51.945 148.265 52.265 ;
        RECT 148.345 51.945 148.665 52.265 ;
        RECT 148.745 51.945 149.065 52.265 ;
        RECT 149.145 51.945 149.465 52.265 ;
        RECT 149.545 51.945 149.865 52.265 ;
        RECT 149.945 51.945 150.265 52.265 ;
        RECT 150.345 51.945 150.665 52.265 ;
        RECT 150.745 51.945 151.065 52.265 ;
        RECT 151.145 51.945 151.465 52.265 ;
        RECT 151.545 51.945 151.865 52.265 ;
        RECT 151.945 51.945 152.265 52.265 ;
        RECT 152.345 51.945 152.665 52.265 ;
        RECT 152.745 51.945 153.065 52.265 ;
        RECT 153.145 51.945 153.465 52.265 ;
        RECT 153.545 51.945 153.865 52.265 ;
        RECT 153.945 51.945 154.265 52.265 ;
        RECT 154.345 51.945 154.665 52.265 ;
        RECT 154.745 51.945 155.065 52.265 ;
        RECT 155.145 51.945 155.465 52.265 ;
        RECT 155.545 51.945 155.865 52.265 ;
        RECT 155.945 51.945 156.265 52.265 ;
        RECT 156.345 51.945 156.665 52.265 ;
        RECT 156.745 51.945 157.065 52.265 ;
        RECT 157.145 51.945 157.465 52.265 ;
        RECT 157.545 51.945 157.865 52.265 ;
        RECT 157.945 51.945 158.265 52.265 ;
        RECT 158.345 51.945 158.665 52.265 ;
        RECT 158.745 51.945 159.065 52.265 ;
        RECT 159.145 51.945 159.465 52.265 ;
        RECT 159.545 51.945 159.865 52.265 ;
        RECT 159.945 51.945 160.265 52.265 ;
        RECT 160.345 51.945 160.665 52.265 ;
        RECT 160.745 51.945 161.065 52.265 ;
        RECT 161.145 51.945 161.465 52.265 ;
        RECT 161.545 51.945 161.865 52.265 ;
        RECT 161.945 51.945 162.265 52.265 ;
        RECT 107.380 44.230 107.700 44.550 ;
        RECT 107.380 43.680 107.700 44.000 ;
      LAYER met4 ;
        RECT -42.900 84.365 161.710 86.090 ;
        RECT -42.900 53.035 -13.290 82.645 ;
        RECT -7.900 53.035 21.710 82.645 ;
        RECT 27.100 53.035 56.710 82.645 ;
        RECT 62.100 53.035 91.710 82.645 ;
        RECT 97.100 53.035 126.710 82.645 ;
        RECT 132.100 53.035 161.710 82.645 ;
        RECT -43.535 51.865 -12.655 52.345 ;
        RECT -8.535 51.865 22.345 52.345 ;
        RECT 26.465 51.865 57.345 52.345 ;
        RECT 61.465 51.865 92.345 52.345 ;
        RECT 96.465 51.865 127.345 52.345 ;
        RECT 131.465 51.865 162.345 52.345 ;
        RECT -43.535 50.905 162.345 51.865 ;
        RECT 107.350 43.650 107.730 50.905 ;
      LAYER via4 ;
        RECT -41.370 84.635 -40.190 85.815 ;
        RECT -39.770 84.635 -38.590 85.815 ;
        RECT -6.370 84.635 -5.190 85.815 ;
        RECT -4.770 84.635 -3.590 85.815 ;
        RECT 28.630 84.635 29.810 85.815 ;
        RECT 30.230 84.635 31.410 85.815 ;
        RECT 63.630 84.635 64.810 85.815 ;
        RECT 65.230 84.635 66.410 85.815 ;
        RECT 98.630 84.635 99.810 85.815 ;
        RECT 100.230 84.635 101.410 85.815 ;
        RECT 133.630 84.635 134.810 85.815 ;
        RECT 135.230 84.635 136.410 85.815 ;
        RECT -41.370 80.885 -40.190 82.065 ;
        RECT -39.770 80.885 -38.590 82.065 ;
        RECT -6.370 80.885 -5.190 82.065 ;
        RECT -4.770 80.885 -3.590 82.065 ;
        RECT 28.630 80.885 29.810 82.065 ;
        RECT 30.230 80.885 31.410 82.065 ;
        RECT 63.630 80.885 64.810 82.065 ;
        RECT 65.230 80.885 66.410 82.065 ;
        RECT 98.630 80.885 99.810 82.065 ;
        RECT 100.230 80.885 101.410 82.065 ;
        RECT 133.630 80.885 134.810 82.065 ;
        RECT 135.230 80.885 136.410 82.065 ;
      LAYER met5 ;
        RECT -41.490 80.765 -38.470 85.935 ;
        RECT -6.490 80.765 -3.470 85.935 ;
        RECT 28.510 80.765 31.530 85.935 ;
        RECT 63.510 80.765 66.530 85.935 ;
        RECT 98.510 80.765 101.530 85.935 ;
        RECT 133.510 80.765 136.530 85.935 ;
  END
END myopamp
END LIBRARY

