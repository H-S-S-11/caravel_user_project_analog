**.subckt analogue_mux_tb
V1 vdd3v3 GND 3.3
V2 VIN1 GND SIN(1.6 1.6 100Meg 0 0)
V3 SEL GND PWL(0 3.3 65n 3.3 70n 0 100n 0)
V4 EN GND PWL(0 0 45n 0 50n 3.3 100n 3.3)
R1 VOUT GND 10k m=1
R2 vdd3v3 VOUT 10k m=1
x2 vdd3v3 VIN0 VOUT VIN1 GND SEL EN analog_mux_2_1
V5 VIN0 GND SIN(1.6 1.6 200Meg 0 0)
**** begin user architecture code


.lib ~/open_sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt


.control
tran 0.1n 100n
plot V(vdd3v3) V(VOUT)
plot V(vdd3v3) VIN0 VIN1 SEL EN
.endc

**** end user architecture code
**.ends

* expanding   symbol:  analog_mux_2_1.sym # of pins=7
* sym_path:
*+ /home/hss11/winhome/skywater-shuttle/caravel_user_project_analog/xschem/analog_mux/analog_mux_2_1.sym
* sch_path:
*+ /home/hss11/winhome/skywater-shuttle/caravel_user_project_analog/xschem/analog_mux/analog_mux_2_1.sch
.subckt analog_mux_2_1  VDD3v3 VIN0 VOUT VIN1 VGND SELECT EN
*.iopin VGND
*.ipin VIN0
*.opin VOUT
*.iopin VDD3v3
*.ipin VIN1
*.ipin EN
*.ipin SELECT
x1 VGND VDD3v3 VIN0 !EN0 EN0 VOUT analogue_switch
x2 VGND VDD3v3 VIN1 !EN1 EN1 VOUT analogue_switch
XM3 !EN1 SELECT VDD3v3 VDD3v3 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM4 !EN1 EN VDD3v3 VDD3v3 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM2 net1 SELECT VGND VGND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM5 !EN1 EN net1 VGND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 EN1 !EN1 VDD3v3 VDD3v3 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM6 EN1 !EN1 VGND VGND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7 !SELECT SELECT VDD3v3 VDD3v3 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM8 !SELECT SELECT VGND VGND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM9 !EN0 EN VDD3v3 VDD3v3 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM10 net2 !SELECT VGND VGND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM11 !EN0 EN net2 VGND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM12 EN0 !EN0 VDD3v3 VDD3v3 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM13 EN0 !EN0 VGND VGND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM14 !EN0 !SELECT VDD3v3 VDD3v3 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  analogue_switch.sym # of pins=6
* sym_path:
*+ /home/hss11/winhome/skywater-shuttle/caravel_user_project_analog/xschem/analog_mux/analogue_switch.sym
* sch_path:
*+ /home/hss11/winhome/skywater-shuttle/caravel_user_project_analog/xschem/analog_mux/analogue_switch.sch
.subckt analogue_switch  VGND VDD3v3 VIN !EN EN VOUT
*.ipin EN
*.ipin VIN
*.opin VOUT
*.ipin !EN
*.iopin VGND
*.iopin VDD3v3
XM2 mid !EN VIN VDD3v3 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM1 VIN EN mid VGND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM3 mid !EN VGND VGND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 VOUT !EN mid VDD3v3 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM5 mid EN VOUT VGND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
.ends

.GLOBAL GND
** flattened .save nodes
.end
