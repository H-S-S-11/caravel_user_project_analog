magic
tech sky130A
magscale 1 2
timestamp 1632865024
<< locali >>
rect 1760 1900 1860 1920
rect 1760 1840 1780 1900
rect 1840 1840 1860 1900
rect 1760 1540 1860 1840
rect 1760 1480 1780 1540
rect 1840 1480 1860 1540
rect 1760 1460 1860 1480
<< viali >>
rect 1780 1840 1840 1900
rect 1780 1480 1840 1540
<< metal1 >>
rect -240 3240 2400 3280
rect -240 3040 2100 3240
rect 2360 3040 2400 3240
rect -240 3000 2400 3040
rect -240 2420 40 3000
rect 480 2720 1620 2760
rect 480 2420 520 2720
rect 820 2420 1620 2720
rect 2060 2460 2400 3000
rect 4560 3000 5600 3200
rect 2720 2720 4420 2760
rect 2720 2600 4080 2720
rect 480 2180 1620 2420
rect 4040 2420 4080 2600
rect 4380 2420 4420 2720
rect 4040 2320 4420 2420
rect 4560 2320 4660 3000
rect 4940 2720 5320 2800
rect 4940 2420 4980 2720
rect 5280 2420 5320 2720
rect 4940 2380 5320 2420
rect 4940 2320 5360 2380
rect 1140 1980 1620 2180
rect -440 1900 1860 1920
rect -440 1840 1780 1900
rect 1840 1840 1860 1900
rect -440 1820 1860 1840
rect 2900 1780 3900 1880
rect 460 1640 2000 1740
rect 460 1420 580 1640
rect 1760 1540 1860 1560
rect 1760 1480 1780 1540
rect 1840 1480 1860 1540
rect 1230 1380 1600 1470
rect -440 1270 540 1350
rect 1500 1340 1600 1380
rect 1760 1340 1860 1480
rect 1500 1240 1860 1340
rect 1900 1320 2000 1640
rect 3800 1280 3900 1780
rect -440 1160 540 1240
rect 460 860 580 1080
rect 1900 860 2000 1220
rect 460 760 2000 860
rect 3800 720 3900 840
rect 2880 620 3900 720
<< via1 >>
rect 2100 3040 2360 3240
rect 520 2420 820 2720
rect 4080 2420 4380 2720
rect 4980 2420 5280 2720
<< metal2 >>
rect 480 2760 840 3400
rect 2060 3240 2400 3400
rect 2060 3040 2100 3240
rect 2360 3040 2400 3240
rect 2060 3000 2400 3040
rect 480 2720 4420 2760
rect 480 2420 520 2720
rect 820 2420 4080 2720
rect 4380 2420 4420 2720
rect 480 2380 4420 2420
rect 4940 2720 5320 3400
rect 4940 2420 4980 2720
rect 5280 2420 5320 2720
rect 4940 2380 5320 2420
use diffamp  diffamp_0
timestamp 1632488633
transform 1 0 4840 0 1 -1080
box -940 980 620 3400
use decision  decision_0
timestamp 1632485541
transform 1 0 2020 0 1 145
box -120 -245 1711 2620
use preamp  preamp_0
timestamp 1632332974
transform 1 0 -145 0 1 115
box -255 -115 1909 2460
<< labels >>
rlabel metal1 -440 1270 -430 1350 1 VP
port 2 n
rlabel metal1 -440 1160 -430 1240 1 VN
port 1 n
rlabel metal1 -440 1820 -420 1920 1 BIASN
port 3 n
rlabel metal1 2060 2760 2400 2800 1 VDD3v3
port 4 n
rlabel metal1 -240 2760 40 2800 1 VDD3v3
port 4 n
rlabel metal2 480 3320 840 3400 1 VGND
port 8 n
rlabel metal2 2060 3320 2400 3400 1 VDD3v3
port 4 n
rlabel metal2 4940 3300 5320 3400 1 VDD1v8
port 9 n
rlabel metal1 5560 3000 5600 3200 1 VOUT
port 10 n
<< end >>
