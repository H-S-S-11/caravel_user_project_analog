magic
tech sky130A
timestamp 1635205324
<< nwell >>
rect 1400 1950 2150 2700
rect 1350 -2650 2150 -2000
<< nnmos >>
rect 980 2470 1050 2520
rect 980 2370 1050 2420
rect 980 2270 1050 2320
rect 980 2140 1050 2190
rect 980 -2240 1050 -2190
rect 980 -2370 1050 -2320
rect 980 -2470 1050 -2420
<< mvpmos >>
rect 1500 2470 1600 2520
rect 1500 2370 1600 2420
rect 1500 2270 1600 2320
rect 1500 2140 1600 2190
rect 1500 -2240 1600 -2190
rect 1500 -2370 1600 -2320
rect 1500 -2470 1600 -2420
<< mvndiff >>
rect 980 2550 1050 2560
rect 980 2530 990 2550
rect 1040 2530 1050 2550
rect 980 2520 1050 2530
rect 980 2460 1050 2470
rect 980 2430 990 2460
rect 1040 2430 1050 2460
rect 980 2420 1050 2430
rect 980 2320 1050 2370
rect 980 2260 1050 2270
rect 980 2200 990 2260
rect 1040 2200 1050 2260
rect 980 2190 1050 2200
rect 980 2130 1050 2140
rect 980 2110 990 2130
rect 1040 2110 1050 2130
rect 980 2100 1050 2110
rect 980 -2160 1050 -2150
rect 980 -2180 990 -2160
rect 1040 -2180 1050 -2160
rect 980 -2190 1050 -2180
rect 980 -2250 1050 -2240
rect 980 -2310 990 -2250
rect 1040 -2310 1050 -2250
rect 980 -2320 1050 -2310
rect 980 -2420 1050 -2370
rect 980 -2480 1050 -2470
rect 980 -2500 990 -2480
rect 1040 -2500 1050 -2480
rect 980 -2510 1050 -2500
<< mvpdiff >>
rect 1500 2550 1600 2560
rect 1500 2530 1510 2550
rect 1590 2530 1600 2550
rect 1500 2520 1600 2530
rect 1500 2460 1600 2470
rect 1500 2430 1510 2460
rect 1590 2430 1600 2460
rect 1500 2420 1600 2430
rect 1500 2360 1600 2370
rect 1500 2330 1510 2360
rect 1590 2330 1600 2360
rect 1500 2320 1600 2330
rect 1500 2260 1600 2270
rect 1500 2200 1510 2260
rect 1590 2200 1600 2260
rect 1500 2190 1600 2200
rect 1500 2130 1600 2140
rect 1500 2110 1510 2130
rect 1590 2110 1600 2130
rect 1500 2100 1600 2110
rect 1500 -2160 1600 -2150
rect 1500 -2180 1510 -2160
rect 1590 -2180 1600 -2160
rect 1500 -2190 1600 -2180
rect 1500 -2250 1600 -2240
rect 1500 -2310 1510 -2250
rect 1590 -2310 1600 -2250
rect 1500 -2320 1600 -2310
rect 1500 -2380 1600 -2370
rect 1500 -2410 1510 -2380
rect 1590 -2410 1600 -2380
rect 1500 -2420 1600 -2410
rect 1500 -2480 1600 -2470
rect 1500 -2500 1510 -2480
rect 1590 -2500 1600 -2480
rect 1500 -2510 1600 -2500
<< mvndiffc >>
rect 990 2530 1040 2550
rect 990 2430 1040 2460
rect 990 2200 1040 2260
rect 990 2110 1040 2130
rect 990 -2180 1040 -2160
rect 990 -2310 1040 -2250
rect 990 -2500 1040 -2480
<< mvpdiffc >>
rect 1510 2530 1590 2550
rect 1510 2430 1590 2460
rect 1510 2330 1590 2360
rect 1510 2200 1590 2260
rect 1510 2110 1590 2130
rect 1510 -2180 1590 -2160
rect 1510 -2310 1590 -2250
rect 1510 -2410 1590 -2380
rect 1510 -2500 1590 -2480
<< mvpsubdiff >>
rect 850 2600 1150 2650
rect 650 2550 900 2600
rect 650 2100 700 2550
rect 850 2100 900 2550
rect 650 2050 900 2100
rect 850 2000 1150 2050
rect 850 -2100 1150 -2050
rect 850 -2150 900 -2100
rect 650 -2200 900 -2150
rect 650 -2500 700 -2200
rect 850 -2500 900 -2200
rect 650 -2550 900 -2500
rect 850 -2600 1150 -2550
<< mvnsubdiff >>
rect 1450 2600 1750 2650
rect 1700 2550 2100 2600
rect 1700 2100 1750 2550
rect 2050 2100 2100 2550
rect 1700 2050 2100 2100
rect 1450 2000 1750 2050
rect 1400 -2100 1700 -2050
rect 1650 -2150 1700 -2100
rect 1650 -2200 2100 -2150
rect 1650 -2500 1700 -2200
rect 1650 -2550 2100 -2500
rect 1400 -2600 1700 -2550
<< mvpsubdiffcont >>
rect 700 2100 850 2550
rect 700 -2500 850 -2200
<< mvnsubdiffcont >>
rect 1750 2100 2050 2550
rect 1700 -2500 2100 -2200
<< poly >>
rect 1310 2520 1380 2530
rect 960 2470 980 2520
rect 1050 2470 1320 2520
rect 1370 2470 1500 2520
rect 1600 2470 1620 2520
rect 1310 2460 1380 2470
rect 1090 2420 1160 2430
rect 960 2370 980 2420
rect 1050 2370 1100 2420
rect 1150 2370 1500 2420
rect 1600 2370 1620 2420
rect 1090 2360 1160 2370
rect 1170 2320 1240 2330
rect 960 2270 980 2320
rect 1050 2270 1180 2320
rect 1230 2270 1500 2320
rect 1600 2270 1620 2320
rect 1170 2260 1240 2270
rect 1220 2191 1340 2200
rect 1220 2190 1231 2191
rect 960 2140 980 2190
rect 1050 2141 1231 2190
rect 1331 2190 1340 2191
rect 1331 2141 1500 2190
rect 1050 2140 1500 2141
rect 1600 2140 1620 2190
rect 1220 2130 1340 2140
rect 1220 -2190 1340 -2180
rect 960 -2240 980 -2190
rect 1050 -2240 1230 -2190
rect 1330 -2240 1500 -2190
rect 1600 -2240 1620 -2190
rect 1220 -2250 1340 -2240
rect 1170 -2320 1240 -2310
rect 960 -2370 980 -2320
rect 1050 -2370 1180 -2320
rect 1230 -2370 1500 -2320
rect 1600 -2370 1620 -2320
rect 1170 -2380 1240 -2370
rect 1310 -2420 1380 -2410
rect 960 -2470 980 -2420
rect 1050 -2470 1320 -2420
rect 1370 -2470 1500 -2420
rect 1600 -2470 1620 -2420
rect 1310 -2480 1380 -2470
<< polycont >>
rect 1320 2470 1370 2520
rect 1100 2370 1150 2420
rect 1180 2270 1230 2320
rect 1231 2141 1331 2191
rect 1230 -2240 1330 -2190
rect 1180 -2370 1230 -2320
rect 1320 -2470 1370 -2420
<< locali >>
rect 650 2550 900 2600
rect 850 2460 900 2550
rect 980 2550 1600 2600
rect 980 2530 990 2550
rect 1040 2530 1050 2550
rect 850 2430 990 2460
rect 1040 2430 1050 2460
rect 1100 2430 1150 2550
rect 1500 2530 1510 2550
rect 1590 2530 1600 2550
rect 1700 2550 2100 2600
rect 1700 2460 1750 2550
rect 1500 2430 1510 2460
rect 1590 2430 1750 2460
rect 850 2130 900 2430
rect 1090 2420 1160 2430
rect 1090 2370 1100 2420
rect 1150 2370 1160 2420
rect 1090 2360 1160 2370
rect 1400 2330 1510 2360
rect 1590 2330 1600 2360
rect 1050 2200 1150 2260
rect 1100 2190 1150 2200
rect 1220 2191 1340 2200
rect 1220 2190 1231 2191
rect 1100 2141 1231 2190
rect 1331 2190 1340 2191
rect 1400 2190 1450 2330
rect 1700 2260 1750 2430
rect 1500 2200 1510 2260
rect 1590 2200 1750 2260
rect 1331 2141 1450 2190
rect 1100 2140 1450 2141
rect 1220 2130 1340 2140
rect 850 2110 990 2130
rect 1040 2110 1050 2130
rect 850 2100 1050 2110
rect 650 2050 900 2100
rect 980 2040 1050 2050
rect 980 1900 1050 1980
rect 1400 1970 1450 2140
rect 1500 2110 1510 2130
rect 1590 2110 1600 2130
rect 1500 2100 1600 2110
rect 1700 2100 1750 2200
rect 1700 2050 2100 2100
rect 1400 1920 1550 1970
rect 800 1850 1050 1900
rect 1500 1900 1550 1920
rect 1500 1850 1750 1900
rect 800 -1950 1050 -1900
rect 980 -2100 1050 -1950
rect 1500 -1950 1750 -1900
rect 1500 -1970 1550 -1950
rect 650 -2200 900 -2150
rect 980 -2160 1050 -2150
rect 980 -2180 990 -2160
rect 1040 -2180 1050 -2160
rect 1400 -2020 1550 -1970
rect 1220 -2190 1340 -2180
rect 1400 -2190 1450 -2020
rect 1500 -2160 1600 -2150
rect 1500 -2180 1510 -2160
rect 1590 -2180 1600 -2160
rect 850 -2250 900 -2200
rect 1100 -2240 1230 -2190
rect 1330 -2240 1450 -2190
rect 850 -2310 990 -2250
rect 1040 -2310 1050 -2250
rect 850 -2500 900 -2310
rect 1100 -2480 1150 -2240
rect 1220 -2250 1340 -2240
rect 1400 -2380 1450 -2240
rect 1650 -2200 2150 -2150
rect 1650 -2250 1700 -2200
rect 1500 -2310 1510 -2250
rect 1590 -2310 1700 -2250
rect 1400 -2410 1510 -2380
rect 1590 -2410 1600 -2380
rect 1650 -2480 1700 -2310
rect 650 -2550 900 -2500
rect 980 -2500 990 -2480
rect 1040 -2500 1150 -2480
rect 980 -2510 1150 -2500
rect 1500 -2500 1510 -2480
rect 1590 -2500 1700 -2480
rect 2100 -2500 2150 -2200
rect 1500 -2510 2150 -2500
rect 1650 -2550 2150 -2510
<< viali >>
rect 650 2100 700 2550
rect 700 2100 850 2550
rect 1310 2520 1380 2530
rect 1310 2470 1320 2520
rect 1320 2470 1370 2520
rect 1370 2470 1380 2520
rect 1310 2460 1380 2470
rect 1170 2320 1240 2330
rect 1170 2270 1180 2320
rect 1180 2270 1230 2320
rect 1230 2270 1240 2320
rect 1170 2260 1240 2270
rect 980 2200 990 2260
rect 990 2200 1040 2260
rect 1040 2200 1050 2260
rect 980 1980 1050 2040
rect 1500 2050 1600 2100
rect 1750 2100 2050 2550
rect 2050 2100 2100 2550
rect 980 -2150 1050 -2100
rect 1500 -2150 1600 -2100
rect 650 -2500 700 -2200
rect 700 -2500 850 -2200
rect 1170 -2320 1240 -2310
rect 1170 -2370 1180 -2320
rect 1180 -2370 1230 -2320
rect 1230 -2370 1240 -2320
rect 1170 -2380 1240 -2370
rect 1310 -2420 1380 -2410
rect 1310 -2470 1320 -2420
rect 1320 -2470 1370 -2420
rect 1370 -2470 1380 -2420
rect 1310 -2480 1380 -2470
rect 1700 -2500 2100 -2200
<< metal1 >>
rect 400 2590 900 2600
rect 400 2110 410 2590
rect 590 2550 900 2590
rect 400 2060 420 2110
rect 590 2100 650 2550
rect 850 2100 900 2550
rect 1700 2590 2350 2600
rect 1700 2550 2160 2590
rect 1300 2530 1390 2540
rect 1300 2460 1310 2530
rect 1380 2460 1390 2530
rect 1300 2450 1390 2460
rect 1160 2330 1250 2340
rect 590 2060 900 2100
rect 400 2050 900 2060
rect 970 2260 1060 2270
rect 970 2200 980 2260
rect 1050 2200 1060 2260
rect 1160 2260 1170 2330
rect 1240 2260 1250 2330
rect 1160 2250 1250 2260
rect 970 2110 1060 2200
rect 970 2100 1610 2110
rect 970 2050 1500 2100
rect 1600 2050 1610 2100
rect 1700 2100 1750 2550
rect 2100 2100 2160 2550
rect 1700 2060 2160 2100
rect 2340 2060 2350 2590
rect 1700 2050 2350 2060
rect 970 2040 1610 2050
rect 970 1980 980 2040
rect 1050 1980 1060 2040
rect 970 1970 1060 1980
rect 2750 1150 3200 1550
rect -50 350 0 750
rect 2800 600 3200 1150
rect 2800 200 3300 600
rect 2800 -350 3200 200
rect 2750 -750 3200 -350
rect -50 -1550 0 -1150
rect 970 -2100 1610 -2090
rect 970 -2150 980 -2100
rect 1050 -2150 1500 -2100
rect 1600 -2150 1610 -2100
rect 400 -2160 900 -2150
rect 970 -2160 1610 -2150
rect 1650 -2160 2350 -2150
rect 400 -2540 410 -2160
rect 590 -2200 900 -2160
rect 590 -2500 650 -2200
rect 850 -2500 900 -2200
rect 1650 -2200 2160 -2160
rect 1160 -2310 1250 -2300
rect 1160 -2380 1170 -2310
rect 1240 -2380 1250 -2310
rect 1160 -2390 1250 -2380
rect 1300 -2410 1390 -2400
rect 1300 -2480 1310 -2410
rect 1380 -2480 1390 -2410
rect 1300 -2490 1390 -2480
rect 590 -2540 900 -2500
rect 400 -2550 900 -2540
rect 1650 -2500 1700 -2200
rect 2100 -2500 2160 -2200
rect 1650 -2540 2160 -2500
rect 2340 -2540 2350 -2160
rect 1650 -2550 2350 -2540
<< via1 >>
rect 410 2110 590 2590
rect 420 2060 590 2110
rect 1310 2460 1380 2530
rect 1170 2260 1240 2330
rect 2160 2060 2340 2590
rect 410 -2540 590 -2160
rect 1170 -2380 1240 -2310
rect 1310 -2480 1380 -2410
rect 2160 -2540 2340 -2160
<< metal2 >>
rect 100 2590 600 2750
rect 100 2110 410 2590
rect 100 2060 420 2110
rect 590 2060 600 2590
rect 100 1850 600 2060
rect 1150 2330 1250 2750
rect 1150 2260 1170 2330
rect 1240 2260 1250 2330
rect 100 -50 600 0
rect 100 -2160 600 -1900
rect 100 -2540 410 -2160
rect 590 -2540 600 -2160
rect 100 -2700 600 -2540
rect 1150 -2310 1250 2260
rect 1150 -2380 1170 -2310
rect 1240 -2380 1250 -2310
rect 1150 -2700 1250 -2380
rect 1300 2530 1400 2750
rect 1300 2460 1310 2530
rect 1380 2460 1400 2530
rect 1300 -2410 1400 2460
rect 2150 2590 2650 2750
rect 2150 2060 2160 2590
rect 2340 2060 2650 2590
rect 2150 1850 2650 2060
rect 2150 -50 2650 0
rect 1300 -2480 1310 -2410
rect 1380 -2480 1400 -2410
rect 1300 -2700 1400 -2480
rect 2150 -2160 2650 -1900
rect 2150 -2540 2160 -2160
rect 2340 -2540 2650 -2160
rect 2150 -2700 2650 -2540
use analog_switch  analog_switch_1
timestamp 1634764606
transform 1 0 500 0 1 -1150
box -500 -750 2250 1100
use analog_switch  analog_switch_0
timestamp 1634764606
transform 1 0 500 0 1 750
box -500 -750 2250 1100
<< labels >>
rlabel locali 990 -2040 1040 -1990 1 EN0
rlabel locali 1450 -2010 1490 -1980 1 ENB0
rlabel locali 990 1910 1040 1960 1 EN1
rlabel locali 1510 1910 1540 1960 1 ENB1
rlabel metal2 100 2700 600 2750 1 VGND
port 1 n
rlabel metal2 2150 2700 2650 2750 1 VPWR
port 2 n
rlabel metal1 -50 350 -20 750 1 VIN1
port 3 n
rlabel metal1 -50 -1550 -20 -1150 1 VIN0
port 4 n
rlabel metal1 3250 200 3300 600 1 VOUT
port 5 n
rlabel metal2 1150 2700 1250 2750 1 EN
port 6 n
rlabel metal2 1150 -2700 1250 -2650 1 EN
port 6 n
rlabel metal2 1300 -2700 1400 -2650 1 SELECT
port 7 n
rlabel metal2 1300 2700 1400 2750 1 SELECT
port 7 n
rlabel locali 1070 2560 1110 2590 1 !SELECT
rlabel metal2 100 -2700 600 -2650 1 VGND
port 1 n
rlabel metal2 2150 -2700 2650 -2650 1 VPWR
port 2 n
<< end >>
