magic
tech sky130A
magscale 1 4
timestamp 1632400215
<< nwell >>
rect -619 -1946 619 1946
<< pmos >>
rect -226 1108 -154 1508
rect -36 1108 36 1508
rect 154 1108 226 1508
rect -226 236 -154 636
rect -36 236 36 636
rect 154 236 226 636
rect -226 -636 -154 -236
rect -36 -636 36 -236
rect 154 -636 226 -236
rect -226 -1508 -154 -1108
rect -36 -1508 36 -1108
rect 154 -1508 226 -1108
<< pdiff >>
rect -343 1484 -226 1508
rect -343 1132 -319 1484
rect -251 1132 -226 1484
rect -343 1108 -226 1132
rect -154 1484 -36 1508
rect -154 1132 -129 1484
rect -61 1132 -36 1484
rect -154 1108 -36 1132
rect 36 1484 154 1508
rect 36 1132 61 1484
rect 129 1132 154 1484
rect 36 1108 154 1132
rect 226 1484 343 1508
rect 226 1132 251 1484
rect 319 1132 343 1484
rect 226 1108 343 1132
rect -343 612 -226 636
rect -343 260 -319 612
rect -251 260 -226 612
rect -343 236 -226 260
rect -154 612 -36 636
rect -154 260 -129 612
rect -61 260 -36 612
rect -154 236 -36 260
rect 36 612 154 636
rect 36 260 61 612
rect 129 260 154 612
rect 36 236 154 260
rect 226 612 343 636
rect 226 260 251 612
rect 319 260 343 612
rect 226 236 343 260
rect -343 -260 -226 -236
rect -343 -612 -319 -260
rect -251 -612 -226 -260
rect -343 -636 -226 -612
rect -154 -260 -36 -236
rect -154 -612 -129 -260
rect -61 -612 -36 -260
rect -154 -636 -36 -612
rect 36 -260 154 -236
rect 36 -612 61 -260
rect 129 -612 154 -260
rect 36 -636 154 -612
rect 226 -260 343 -236
rect 226 -612 251 -260
rect 319 -612 343 -260
rect 226 -636 343 -612
rect -343 -1132 -226 -1108
rect -343 -1484 -319 -1132
rect -251 -1484 -226 -1132
rect -343 -1508 -226 -1484
rect -154 -1132 -36 -1108
rect -154 -1484 -129 -1132
rect -61 -1484 -36 -1132
rect -154 -1508 -36 -1484
rect 36 -1132 154 -1108
rect 36 -1484 61 -1132
rect 129 -1484 154 -1132
rect 36 -1508 154 -1484
rect 226 -1132 343 -1108
rect 226 -1484 251 -1132
rect 319 -1484 343 -1132
rect 226 -1508 343 -1484
<< pdiffc >>
rect -319 1132 -251 1484
rect -129 1132 -61 1484
rect 61 1132 129 1484
rect 251 1132 319 1484
rect -319 260 -251 612
rect -129 260 -61 612
rect 61 260 129 612
rect 251 260 319 612
rect -319 -612 -251 -260
rect -129 -612 -61 -260
rect 61 -612 129 -260
rect 251 -612 319 -260
rect -319 -1484 -251 -1132
rect -129 -1484 -61 -1132
rect 61 -1484 129 -1132
rect 251 -1484 319 -1132
<< nsubdiff >>
rect -547 1806 -355 1874
rect 355 1806 547 1874
rect -547 1682 -479 1806
rect 479 1682 547 1806
rect -547 -1806 -479 -1682
rect 479 -1806 547 -1682
rect -547 -1874 -355 -1806
rect 355 -1874 547 -1806
<< nsubdiffcont >>
rect -355 1806 355 1874
rect -547 -1682 -479 1682
rect 479 -1682 547 1682
rect -355 -1874 355 -1806
<< poly >>
rect -256 1670 -124 1702
rect -256 1602 -224 1670
rect -156 1602 -124 1670
rect -256 1570 -124 1602
rect 124 1670 256 1702
rect 124 1602 156 1670
rect 224 1602 256 1670
rect 124 1570 256 1602
rect -226 1508 -154 1570
rect -36 1508 36 1560
rect 154 1508 226 1570
rect -226 1056 -154 1108
rect -36 1046 36 1108
rect 154 1056 226 1108
rect -66 1014 66 1046
rect -66 946 -34 1014
rect 34 946 66 1014
rect -66 920 66 946
rect -226 636 -154 700
rect -36 636 36 700
rect 154 636 226 700
rect -226 180 -154 236
rect -36 180 36 236
rect 154 180 226 236
rect -226 -180 227 180
rect -226 -236 -154 -180
rect -36 -236 36 -180
rect 154 -236 226 -180
rect -226 -700 -154 -636
rect -36 -700 36 -636
rect 154 -700 226 -636
rect -226 -730 226 -700
rect -226 -798 -34 -730
rect 34 -798 226 -730
rect -226 -820 226 -798
rect -66 -946 66 -914
rect -66 -1014 -34 -946
rect 34 -1014 66 -946
rect -66 -1046 66 -1014
rect -226 -1108 -154 -1056
rect -36 -1108 36 -1046
rect 154 -1108 226 -1056
rect -226 -1570 -154 -1508
rect -36 -1560 36 -1508
rect 154 -1570 226 -1508
rect -256 -1602 -124 -1570
rect -256 -1670 -224 -1602
rect -156 -1670 -124 -1602
rect -256 -1702 -124 -1670
rect 124 -1602 256 -1570
rect 124 -1670 156 -1602
rect 224 -1670 256 -1602
rect 124 -1702 256 -1670
<< polycont >>
rect -224 1602 -156 1670
rect 156 1602 224 1670
rect -34 946 34 1014
rect -34 -798 34 -730
rect -34 -1014 34 -946
rect -224 -1670 -156 -1602
rect 156 -1670 224 -1602
<< locali >>
rect -547 1806 -355 1874
rect 355 1806 547 1874
rect -547 1682 -479 1806
rect 479 1682 547 1806
rect -256 1602 -224 1670
rect -156 1602 -124 1670
rect 124 1602 156 1670
rect 224 1602 256 1670
rect -319 1484 -251 1516
rect -319 1100 -251 1132
rect -129 1484 -61 1516
rect -129 1100 -61 1132
rect 61 1484 129 1516
rect 61 1100 129 1132
rect 251 1484 319 1516
rect 251 1100 319 1132
rect -66 946 -34 1014
rect 34 946 66 1014
rect -319 612 -251 644
rect -319 228 -251 260
rect -129 612 -61 644
rect -129 228 -61 260
rect 61 612 129 644
rect 61 228 129 260
rect 251 612 319 644
rect 251 228 319 260
rect -319 -260 -251 -228
rect -319 -644 -251 -612
rect -129 -260 -61 -228
rect -129 -644 -61 -612
rect 61 -260 129 -228
rect 61 -644 129 -612
rect 251 -260 319 -228
rect 251 -644 319 -612
rect -66 -798 -34 -730
rect 34 -798 66 -730
rect -66 -1014 -34 -946
rect 34 -1014 66 -946
rect -319 -1132 -251 -1100
rect -319 -1516 -251 -1484
rect -129 -1132 -61 -1100
rect -129 -1516 -61 -1484
rect 61 -1132 129 -1100
rect 61 -1516 129 -1484
rect 251 -1132 319 -1100
rect 251 -1516 319 -1484
rect -256 -1670 -224 -1602
rect -156 -1670 -124 -1602
rect 124 -1670 156 -1602
rect 224 -1670 256 -1602
rect -547 -1806 -479 -1682
rect 479 -1806 547 -1682
rect -547 -1874 -355 -1806
rect 355 -1874 547 -1806
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -513 -1840 513 1840
string parameters w 1 l 0.18 m 4 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
