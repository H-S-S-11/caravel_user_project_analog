magic
tech sky130A
magscale 1 10000
timestamp 1632485541
<< nwell >>
rect 1718137 3700000 1850000 5200000
<< pwell >>
rect 3500000 4800000 3800000 5300000
rect 3500000 3500000 4300000 3550000
rect 3500000 1800000 3900000 3400000
<< locali >>
rect 3200000 12400000 3600000 12500000
rect 5100000 12400000 5450000 12500000
rect 300000 11600000 1800000 11700000
rect 50000 9050000 2100000 11550000
rect 3200000 10300000 5450000 12400000
rect 2050000 9000000 2100000 9050000
rect 3500000 9400000 4300000 9800000
rect 6000000 9250000 6400000 9350000
rect 7900000 9250000 8200000 9350000
rect 3500000 8050000 4300000 8500000
rect 50000 6700000 650000 7550000
rect 3500000 6350000 3800000 8050000
rect 4800000 6650000 5150000 9250000
rect 6000000 7150000 8200000 9250000
rect 500000 5950000 1350000 6150000
rect 300000 5900000 1350000 5950000
rect 3500000 6000000 4600000 6100000
rect 3500000 5900000 4500000 6000000
rect 300000 5600000 1350000 5650000
rect 500000 5400000 1350000 5600000
rect 3500000 5300000 3700000 5900000
rect 50000 4050000 650000 4900000
rect 3500000 3550000 3800000 5300000
rect 4800000 4950000 4850000 6650000
rect 7500000 5300000 8250000 6300000
rect 3500000 3100000 4300000 3550000
rect 50000 0 2100000 2550000
rect 4800000 2900000 5150000 4950000
rect 4750000 2300000 5150000 2900000
rect 6050000 2250000 8250000 4450000
rect 3500000 1800000 4300000 2200000
rect 3200000 -900000 5450000 1300000
<< viali >>
rect 3600000 12400000 5100000 12900000
rect 300000 11700000 1800000 12200000
rect 3500000 8500000 4300000 9400000
rect 6400000 9250000 7900000 9750000
rect 1350000 6350000 1850000 7900000
rect 300000 5950000 500000 6150000
rect 300000 5400000 500000 5600000
rect 4150000 5400000 4450000 5700000
rect 1400000 3700000 1850000 5200000
rect 4850000 4950000 5150000 6650000
rect 6350000 4950000 7150000 6650000
rect 3500000 2200000 4300000 3100000
<< metal1 >>
rect 200000 12200000 1900000 13100000
rect 3500000 12900000 8000000 13100000
rect 3500000 12400000 3600000 12900000
rect 5100000 12400000 8000000 12900000
rect 3500000 12300000 8000000 12400000
rect 200000 11700000 300000 12200000
rect 1800000 11700000 1900000 12200000
rect 200000 11600000 1900000 11700000
rect 6300000 9750000 8000000 12300000
rect 3400000 9400000 4550000 9500000
rect 3400000 9300000 3500000 9400000
rect 1250000 8600000 3500000 9300000
rect 1250000 7900000 1950000 8600000
rect 3400000 8500000 3500000 8600000
rect 4300000 8500000 4550000 9400000
rect 6300000 9250000 6400000 9750000
rect 7900000 9250000 8000000 9750000
rect 6300000 9150000 8000000 9250000
rect 3400000 8400000 4550000 8500000
rect 1250000 6350000 1350000 7900000
rect 1850000 6350000 1950000 7900000
rect 1250000 6250000 1950000 6350000
rect -600000 6150000 600000 6250000
rect -600000 5950000 300000 6150000
rect 500000 5950000 600000 6150000
rect -600000 5850000 600000 5950000
rect 4050000 5700000 4550000 8400000
rect -600000 5600000 600000 5700000
rect -600000 5400000 300000 5600000
rect 500000 5400000 600000 5600000
rect -600000 5300000 600000 5400000
rect 4050000 5400000 4150000 5700000
rect 4450000 5400000 4550000 5700000
rect 4050000 5300000 4550000 5400000
rect 4750000 6650000 7250000 6750000
rect 1250000 5200000 1950000 5300000
rect 1250000 3700000 1400000 5200000
rect 1850000 3700000 1950000 5200000
rect 4750000 4950000 4850000 6650000
rect 5150000 4950000 6350000 6650000
rect 7150000 4950000 7250000 6650000
rect 4750000 4850000 7250000 4950000
rect 1250000 3000000 1950000 3700000
rect 3400000 3100000 4400000 3200000
rect 3400000 3000000 3500000 3100000
rect 1250000 2300000 3500000 3000000
rect 3350000 2200000 3500000 2300000
rect 4300000 2200000 4400000 3100000
rect 3350000 2100000 4400000 2200000
use sky130_fd_pr__pfet_g5v0d10v5_CABTE7  sky130_fd_pr__pfet_g5v0d10v5_CABTE7_0
timestamp 1632332974
transform 1 0 1065000 0 1 5780000
box -1540000 -6255000 1540000 6255000
use sky130_fd_pr__nfet_03v3_nvt_BKHJCF  sky130_fd_pr__nfet_03v3_nvt_BKHJCF_0
timestamp 1632337456
transform 1 0 4315000 0 1 5790000
box -1440000 -7015000 1440000 7015000
use sky130_fd_pr__nfet_03v3_nvt_NAHJCF  sky130_fd_pr__nfet_03v3_nvt_NAHJCF_0
timestamp 1632334879
transform 1 0 7115000 0 1 5805000
box -1440000 -3880000 1440000 3880000
<< labels >>
rlabel metal1 200000 12900000 1900000 13100000 1 VPWR
rlabel metal1 1250000 6250000 1950000 8000000 1 VOP
rlabel metal1 1250000 3600000 1950000 5300000 1 VON
rlabel metal1 -600000 5850000 -500000 6250000 1 VPAMP
rlabel metal1 -600000 5300000 -500000 5700000 1 VNAMP
rlabel metal1 6250000 4850000 7250000 6750000 1 ISINK
rlabel metal1 3500000 12900000 8000000 13100000 1 VGND
<< end >>
