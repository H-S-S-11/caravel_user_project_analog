magic
tech sky130A
magscale 1 2
timestamp 1632337456
<< nwell >>
rect 60 1720 270 1770
rect 60 1190 270 1230
rect 40 1180 270 1190
rect 40 1170 120 1180
rect 40 1130 120 1140
rect 40 1110 270 1130
rect 40 1060 120 1110
rect 280 740 370 1040
<< pwell >>
rect 700 960 760 1060
rect 700 700 860 710
rect 700 360 780 680
<< locali >>
rect 640 2480 720 2500
rect 1020 2480 1090 2500
rect 60 2320 360 2340
rect 10 1810 420 2310
rect 640 2060 1090 2480
rect 410 1800 420 1810
rect 700 1880 860 1960
rect 1200 1850 1280 1870
rect 1580 1850 1640 1870
rect 700 1610 860 1700
rect 10 1340 130 1510
rect 700 1270 760 1610
rect 960 1330 1030 1850
rect 1200 1430 1640 1850
rect 100 1190 270 1230
rect 60 1180 270 1190
rect 700 1200 920 1220
rect 700 1180 900 1200
rect 60 1120 270 1130
rect 100 1080 270 1120
rect 700 1060 740 1180
rect 10 810 130 980
rect 700 710 760 1060
rect 960 990 970 1330
rect 1500 1060 1650 1260
rect 700 620 860 710
rect 10 0 420 510
rect 960 580 1030 990
rect 950 460 1030 580
rect 1210 450 1650 890
rect 700 360 860 440
rect 640 -180 1090 260
<< viali >>
rect 720 2480 1020 2580
rect 60 2340 360 2440
rect 700 1700 860 1880
rect 1280 1850 1580 1950
rect 270 1270 370 1580
rect 60 1190 100 1230
rect 60 1080 100 1120
rect 830 1080 890 1140
rect 280 740 370 1040
rect 970 990 1030 1330
rect 1270 990 1430 1330
rect 700 440 860 620
<< metal1 >>
rect 40 2440 380 2620
rect 700 2580 1600 2620
rect 700 2480 720 2580
rect 1020 2480 1600 2580
rect 700 2460 1600 2480
rect 40 2340 60 2440
rect 360 2340 380 2440
rect 40 2320 380 2340
rect 1260 1950 1600 2460
rect 680 1880 910 1900
rect 680 1860 700 1880
rect 250 1720 700 1860
rect 250 1580 390 1720
rect 680 1700 700 1720
rect 860 1700 910 1880
rect 1260 1850 1280 1950
rect 1580 1850 1600 1950
rect 1260 1830 1600 1850
rect 680 1680 910 1700
rect 250 1270 270 1580
rect 370 1270 390 1580
rect 250 1250 390 1270
rect -120 1230 120 1250
rect -120 1190 60 1230
rect 100 1190 120 1230
rect -120 1170 120 1190
rect 810 1140 910 1680
rect -120 1120 120 1140
rect -120 1080 60 1120
rect 100 1080 120 1120
rect -120 1060 120 1080
rect 810 1080 830 1140
rect 890 1080 910 1140
rect 810 1060 910 1080
rect 950 1330 1450 1350
rect 250 1040 390 1060
rect 250 740 280 1040
rect 370 740 390 1040
rect 950 990 970 1330
rect 1030 990 1270 1330
rect 1430 990 1450 1330
rect 950 970 1450 990
rect 250 600 390 740
rect 680 620 880 640
rect 680 600 700 620
rect 250 460 700 600
rect 670 440 700 460
rect 860 440 880 620
rect 670 420 880 440
use sky130_fd_pr__nfet_03v3_nvt_NAHJCF  sky130_fd_pr__nfet_03v3_nvt_NAHJCF_0
timestamp 1632334879
transform 1 0 1423 0 1 1161
box -288 -776 288 776
use sky130_fd_pr__nfet_03v3_nvt_BKHJCF  sky130_fd_pr__nfet_03v3_nvt_BKHJCF_0
timestamp 1632337456
transform 1 0 863 0 1 1158
box -288 -1403 288 1403
use sky130_fd_pr__pfet_g5v0d10v5_CABTE7  sky130_fd_pr__pfet_g5v0d10v5_CABTE7_0
timestamp 1632332974
transform 1 0 213 0 1 1156
box -308 -1251 308 1251
<< labels >>
rlabel metal1 40 2580 380 2620 1 VPWR
rlabel metal1 250 1250 390 1600 1 VOP
rlabel metal1 250 720 390 1060 1 VON
rlabel metal1 -120 1170 -100 1250 1 VPAMP
rlabel metal1 -120 1060 -100 1140 1 VNAMP
rlabel metal1 1250 970 1450 1350 1 ISINK
rlabel metal1 700 2580 1600 2620 1 VGND
<< end >>
