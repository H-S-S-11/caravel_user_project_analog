**.subckt analogue_switch_tb
x1 VIN GND vdd3v3 ENB EN VOUT analogue_switch
V1 vdd3v3 GND 3.3
V2 VIN GND SIN(1.6 1.6 100Meg 0 0)
V3 ENB GND PWL(0 3.3 45n 3.3 50n 0 100n 0)
V4 EN GND PWL(0 0 45n 0 50n 3.3 100n 3.3)
R1 VOUT GND 10k m=1
R2 vdd3v3 VOUT 10k m=1
**** begin user architecture code


.lib ~/open_sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt


.control
tran 0.1n 100n
plot V(vdd3v3) V(VOUT) VIN ENB EN
plot I(V1) I(V2) I(R1)
.endc

**** end user architecture code
**.ends

* expanding   symbol:  analogue_switch.sym # of pins=6
* sym_path: /home/hss11/winhome/caravel_user_project_analog/xschem/analogue_switch.sym
* sch_path: /home/hss11/winhome/caravel_user_project_analog/xschem/analogue_switch.sch
.subckt analogue_switch  VIN VGND VDD3v3 !EN EN VOUT
*.iopin VGND
*.iopin VDD3v3
*.ipin EN
*.ipin VIN
*.ipin !EN
*.opin VOUT
XM2 VOUT !EN VIN VDD3v3 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=15 m=15 
XM1 VIN EN VOUT VGND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10 
.ends

.GLOBAL GND
** flattened .save nodes
.end
