magic
tech sky130A
magscale 1 2
timestamp 1635946216
<< pwell >>
rect -284 -126 284 126
<< mvnmos >>
rect -200 -100 200 100
<< mvndiff >>
rect -258 85 -200 100
rect -258 51 -246 85
rect -212 51 -200 85
rect -258 17 -200 51
rect -258 -17 -246 17
rect -212 -17 -200 17
rect -258 -51 -200 -17
rect -258 -85 -246 -51
rect -212 -85 -200 -51
rect -258 -100 -200 -85
rect 200 85 258 100
rect 200 51 212 85
rect 246 51 258 85
rect 200 17 258 51
rect 200 -17 212 17
rect 246 -17 258 17
rect 200 -51 258 -17
rect 200 -85 212 -51
rect 246 -85 258 -51
rect 200 -100 258 -85
<< mvndiffc >>
rect -246 51 -212 85
rect -246 -17 -212 17
rect -246 -85 -212 -51
rect 212 51 246 85
rect 212 -17 246 17
rect 212 -85 246 -51
<< poly >>
rect -200 172 200 188
rect -200 138 -153 172
rect -119 138 -85 172
rect -51 138 -17 172
rect 17 138 51 172
rect 85 138 119 172
rect 153 138 200 172
rect -200 100 200 138
rect -200 -138 200 -100
rect -200 -172 -153 -138
rect -119 -172 -85 -138
rect -51 -172 -17 -138
rect 17 -172 51 -138
rect 85 -172 119 -138
rect 153 -172 200 -138
rect -200 -188 200 -172
<< polycont >>
rect -153 138 -119 172
rect -85 138 -51 172
rect -17 138 17 172
rect 51 138 85 172
rect 119 138 153 172
rect -153 -172 -119 -138
rect -85 -172 -51 -138
rect -17 -172 17 -138
rect 51 -172 85 -138
rect 119 -172 153 -138
<< locali >>
rect -200 138 -161 172
rect -119 138 -89 172
rect -51 138 -17 172
rect 17 138 51 172
rect 89 138 119 172
rect 161 138 200 172
rect -246 85 -212 104
rect -246 17 -212 19
rect -246 -19 -212 -17
rect -246 -104 -212 -85
rect 212 85 246 104
rect 212 17 246 19
rect 212 -19 246 -17
rect 212 -104 246 -85
rect -200 -172 -161 -138
rect -119 -172 -89 -138
rect -51 -172 -17 -138
rect 17 -172 51 -138
rect 89 -172 119 -138
rect 161 -172 200 -138
<< viali >>
rect -161 138 -153 172
rect -153 138 -127 172
rect -89 138 -85 172
rect -85 138 -55 172
rect -17 138 17 172
rect 55 138 85 172
rect 85 138 89 172
rect 127 138 153 172
rect 153 138 161 172
rect -246 51 -212 53
rect -246 19 -212 51
rect -246 -51 -212 -19
rect -246 -53 -212 -51
rect 212 51 246 53
rect 212 19 246 51
rect 212 -51 246 -19
rect 212 -53 246 -51
rect -161 -172 -153 -138
rect -153 -172 -127 -138
rect -89 -172 -85 -138
rect -85 -172 -55 -138
rect -17 -172 17 -138
rect 55 -172 85 -138
rect 85 -172 89 -138
rect 127 -172 153 -138
rect 153 -172 161 -138
<< metal1 >>
rect -196 172 196 178
rect -196 138 -161 172
rect -127 138 -89 172
rect -55 138 -17 172
rect 17 138 55 172
rect 89 138 127 172
rect 161 138 196 172
rect -196 132 196 138
rect -252 53 -206 100
rect -252 19 -246 53
rect -212 19 -206 53
rect -252 -19 -206 19
rect -252 -53 -246 -19
rect -212 -53 -206 -19
rect -252 -100 -206 -53
rect 206 53 252 100
rect 206 19 212 53
rect 246 19 252 53
rect 206 -19 252 19
rect 206 -53 212 -19
rect 246 -53 252 -19
rect 206 -100 252 -53
rect -196 -138 196 -132
rect -196 -172 -161 -138
rect -127 -172 -89 -138
rect -55 -172 -17 -138
rect 17 -172 55 -138
rect 89 -172 127 -138
rect 161 -172 196 -138
rect -196 -178 196 -172
<< end >>
