magic
tech sky130A
magscale 1 2
timestamp 1635946216
<< error_s >>
rect 2117 8670 2323 8804
rect 3117 8670 3323 8804
rect 1900 8043 1930 8575
rect 1966 8109 1996 8509
rect 2452 8109 2482 8509
rect 2518 8043 2548 8575
rect 2900 8043 2930 8575
rect 2966 8109 2996 8509
rect 3452 8109 3482 8509
rect 3518 8043 3548 8575
rect 1900 7303 1930 7835
rect 1966 7369 1996 7769
rect 2452 7369 2482 7769
rect 2518 7303 2548 7835
rect 2900 7303 2930 7835
rect 2966 7369 2996 7769
rect 3452 7369 3482 7769
rect 3518 7303 3548 7835
rect 2114 7065 2320 7199
rect 3114 7065 3320 7199
rect 11835 7010 12041 7144
rect 12735 7010 12941 7144
rect 13635 7010 13841 7144
rect 14535 7010 14741 7144
rect 15435 7010 15587 7144
rect 11618 6383 11648 6915
rect 11684 6449 11714 6849
rect 12170 6449 12200 6849
rect 12236 6383 12266 6915
rect 12518 6383 12548 6915
rect 12584 6449 12614 6849
rect 13070 6449 13100 6849
rect 13136 6383 13166 6915
rect 13418 6383 13448 6915
rect 13484 6449 13514 6849
rect 13970 6449 14000 6849
rect 14036 6383 14066 6915
rect 14318 6383 14327 6915
rect -1346 5949 -1186 5985
rect -1222 5867 -1186 5949
rect -1346 5831 -1186 5867
rect -712 5949 -486 5985
rect -712 5867 -676 5949
rect -522 5867 -486 5949
rect -712 5831 -486 5867
rect -12 5949 214 5985
rect -12 5867 24 5949
rect 178 5867 214 5949
rect -12 5831 214 5867
rect 688 5949 914 5985
rect 688 5867 724 5949
rect 878 5867 914 5949
rect 688 5831 914 5867
rect 1388 5949 1614 5985
rect 1388 5867 1424 5949
rect 1578 5867 1614 5949
rect 1388 5831 1614 5867
rect 2088 5949 2314 5985
rect 2088 5867 2124 5949
rect 2278 5867 2314 5949
rect 2088 5831 2314 5867
rect 3788 5949 4014 5985
rect 3788 5867 3824 5949
rect 3978 5867 4014 5949
rect 3788 5831 4014 5867
rect 4488 5949 4714 5985
rect 4488 5867 4524 5949
rect 4678 5867 4714 5949
rect 4488 5831 4714 5867
rect 5188 5949 5414 5985
rect 5188 5867 5224 5949
rect 5378 5867 5414 5949
rect 5188 5831 5414 5867
rect 5888 5949 6114 5985
rect 5888 5867 5924 5949
rect 6078 5867 6114 5949
rect 5888 5831 6114 5867
rect 6588 5949 6814 5985
rect 6588 5867 6624 5949
rect 6778 5867 6814 5949
rect 6588 5831 6814 5867
rect 7288 5949 7514 5985
rect 7288 5867 7324 5949
rect 7478 5867 7514 5949
rect 7288 5831 7514 5867
rect 7988 5949 8214 5985
rect 7988 5867 8024 5949
rect 8178 5867 8214 5949
rect 7988 5831 8214 5867
rect 8688 5949 8914 5985
rect 8688 5867 8724 5949
rect 8878 5867 8914 5949
rect 8688 5831 8914 5867
rect 9388 5949 9614 5985
rect 9388 5867 9424 5949
rect 9578 5867 9614 5949
rect 9388 5831 9614 5867
rect 10088 5949 10314 5985
rect 10088 5867 10124 5949
rect 10278 5867 10314 5949
rect 10088 5831 10314 5867
rect -1328 5668 -1326 5702
rect -1292 5668 -1288 5702
rect -628 5668 -626 5702
rect -592 5668 -588 5702
rect 72 5668 74 5702
rect 108 5668 112 5702
rect 772 5668 774 5702
rect 808 5668 812 5702
rect 1472 5668 1474 5702
rect 1508 5668 1512 5702
rect 2172 5668 2174 5702
rect 2208 5668 2212 5702
rect 3872 5668 3874 5702
rect 3908 5668 3912 5702
rect 4572 5668 4574 5702
rect 4608 5668 4612 5702
rect 5272 5668 5274 5702
rect 5308 5668 5312 5702
rect 5972 5668 5974 5702
rect 6008 5668 6012 5702
rect 6672 5668 6674 5702
rect 6708 5668 6712 5702
rect 7372 5668 7374 5702
rect 7408 5668 7412 5702
rect 8072 5668 8074 5702
rect 8108 5668 8112 5702
rect 8772 5668 8774 5702
rect 8808 5668 8812 5702
rect 9472 5668 9474 5702
rect 9508 5668 9512 5702
rect 10172 5668 10174 5702
rect 10208 5668 10212 5702
rect 11618 5643 11648 6175
rect 11684 5709 11714 6109
rect 12170 5709 12200 6109
rect 12236 5643 12266 6175
rect 12518 5643 12548 6175
rect 12584 5709 12614 6109
rect 13070 5709 13100 6109
rect 13136 5643 13166 6175
rect 13418 5643 13448 6175
rect 13484 5709 13514 6109
rect 13970 5709 14000 6109
rect 14036 5643 14066 6175
rect 14318 5643 14327 6175
rect -1196 5564 -1162 5566
rect -754 5564 -720 5566
rect -496 5564 -462 5566
rect -54 5564 -20 5566
rect 204 5564 238 5566
rect 646 5564 680 5566
rect 904 5564 938 5566
rect 1346 5564 1380 5566
rect 1604 5564 1638 5566
rect 2046 5564 2080 5566
rect 2304 5564 2338 5566
rect 3746 5564 3780 5566
rect 4004 5564 4038 5566
rect 4446 5564 4480 5566
rect 4704 5564 4738 5566
rect 5146 5564 5180 5566
rect 5404 5564 5438 5566
rect 5846 5564 5880 5566
rect 6104 5564 6138 5566
rect 6546 5564 6580 5566
rect 6804 5564 6838 5566
rect 7246 5564 7280 5566
rect 7504 5564 7538 5566
rect 7946 5564 7980 5566
rect 8204 5564 8238 5566
rect 8646 5564 8680 5566
rect 8904 5564 8938 5566
rect 9346 5564 9380 5566
rect 9604 5564 9638 5566
rect 10046 5564 10080 5566
rect 10304 5564 10338 5566
rect -1196 5548 -1162 5550
rect -754 5548 -720 5550
rect -496 5548 -462 5550
rect -54 5548 -20 5550
rect 204 5548 238 5550
rect 646 5548 680 5550
rect 904 5548 938 5550
rect 1346 5548 1380 5550
rect 1604 5548 1638 5550
rect 2046 5548 2080 5550
rect 2304 5548 2338 5550
rect 3746 5548 3780 5550
rect 4004 5548 4038 5550
rect 4446 5548 4480 5550
rect 4704 5548 4738 5550
rect 5146 5548 5180 5550
rect 5404 5548 5438 5550
rect 5846 5548 5880 5550
rect 6104 5548 6138 5550
rect 6546 5548 6580 5550
rect 6804 5548 6838 5550
rect 7246 5548 7280 5550
rect 7504 5548 7538 5550
rect 7946 5548 7980 5550
rect 8204 5548 8238 5550
rect 8646 5548 8680 5550
rect 8904 5548 8938 5550
rect 9346 5548 9380 5550
rect 9604 5548 9638 5550
rect 10046 5548 10080 5550
rect 10304 5548 10338 5550
rect -1196 5510 -1162 5512
rect -754 5510 -720 5512
rect -496 5510 -462 5512
rect -54 5510 -20 5512
rect 204 5510 238 5512
rect 646 5510 680 5512
rect 904 5510 938 5512
rect 1346 5510 1380 5512
rect 1604 5510 1638 5512
rect 2046 5510 2080 5512
rect 2304 5510 2338 5512
rect 3746 5510 3780 5512
rect 4004 5510 4038 5512
rect 4446 5510 4480 5512
rect 4704 5510 4738 5512
rect 5146 5510 5180 5512
rect 5404 5510 5438 5512
rect 5846 5510 5880 5512
rect 6104 5510 6138 5512
rect 6546 5510 6580 5512
rect 6804 5510 6838 5512
rect 7246 5510 7280 5512
rect 7504 5510 7538 5512
rect 7946 5510 7980 5512
rect 8204 5510 8238 5512
rect 8646 5510 8680 5512
rect 8904 5510 8938 5512
rect 9346 5510 9380 5512
rect 9604 5510 9638 5512
rect 10046 5510 10080 5512
rect 10304 5510 10338 5512
rect -1196 5496 -1162 5498
rect -754 5496 -720 5498
rect -496 5496 -462 5498
rect -54 5496 -20 5498
rect 204 5496 238 5498
rect 646 5496 680 5498
rect 904 5496 938 5498
rect 1346 5496 1380 5498
rect 1604 5496 1638 5498
rect 2046 5496 2080 5498
rect 2304 5496 2338 5498
rect 3746 5496 3780 5498
rect 4004 5496 4038 5498
rect 4446 5496 4480 5498
rect 4704 5496 4738 5498
rect 5146 5496 5180 5498
rect 5404 5496 5438 5498
rect 5846 5496 5880 5498
rect 6104 5496 6138 5498
rect 6546 5496 6580 5498
rect 6804 5496 6838 5498
rect 7246 5496 7280 5498
rect 7504 5496 7538 5498
rect 7946 5496 7980 5498
rect 8204 5496 8238 5498
rect 8646 5496 8680 5498
rect 8904 5496 8938 5498
rect 9346 5496 9380 5498
rect 9604 5496 9638 5498
rect 10046 5496 10080 5498
rect 10304 5496 10338 5498
rect -1196 5476 -1162 5478
rect -754 5476 -720 5478
rect -496 5476 -462 5478
rect -54 5476 -20 5478
rect 204 5476 238 5478
rect 646 5476 680 5478
rect 904 5476 938 5478
rect 1346 5476 1380 5478
rect 1604 5476 1638 5478
rect 2046 5476 2080 5478
rect 2304 5476 2338 5478
rect 3746 5476 3780 5478
rect 4004 5476 4038 5478
rect 4446 5476 4480 5478
rect 4704 5476 4738 5478
rect 5146 5476 5180 5478
rect 5404 5476 5438 5478
rect 5846 5476 5880 5478
rect 6104 5476 6138 5478
rect 6546 5476 6580 5478
rect 6804 5476 6838 5478
rect 7246 5476 7280 5478
rect 7504 5476 7538 5478
rect 7946 5476 7980 5478
rect 8204 5476 8238 5478
rect 8646 5476 8680 5478
rect 8904 5476 8938 5478
rect 9346 5476 9380 5478
rect 9604 5476 9638 5478
rect 10046 5476 10080 5478
rect 10304 5476 10338 5478
rect -1196 5438 -1162 5440
rect -754 5438 -720 5440
rect -496 5438 -462 5440
rect -54 5438 -20 5440
rect 204 5438 238 5440
rect 646 5438 680 5440
rect 904 5438 938 5440
rect 1346 5438 1380 5440
rect 1604 5438 1638 5440
rect 2046 5438 2080 5440
rect 2304 5438 2338 5440
rect 3746 5438 3780 5440
rect 4004 5438 4038 5440
rect 4446 5438 4480 5440
rect 4704 5438 4738 5440
rect 5146 5438 5180 5440
rect 5404 5438 5438 5440
rect 5846 5438 5880 5440
rect 6104 5438 6138 5440
rect 6546 5438 6580 5440
rect 6804 5438 6838 5440
rect 7246 5438 7280 5440
rect 7504 5438 7538 5440
rect 7946 5438 7980 5440
rect 8204 5438 8238 5440
rect 8646 5438 8680 5440
rect 8904 5438 8938 5440
rect 9346 5438 9380 5440
rect 9604 5438 9638 5440
rect 10046 5438 10080 5440
rect 10304 5438 10338 5440
rect -1196 5428 -1162 5430
rect -754 5428 -720 5430
rect -496 5428 -462 5430
rect -54 5428 -20 5430
rect 204 5428 238 5430
rect 646 5428 680 5430
rect 904 5428 938 5430
rect 1346 5428 1380 5430
rect 1604 5428 1638 5430
rect 2046 5428 2080 5430
rect 2304 5428 2338 5430
rect 3746 5428 3780 5430
rect 4004 5428 4038 5430
rect 4446 5428 4480 5430
rect 4704 5428 4738 5430
rect 5146 5428 5180 5430
rect 5404 5428 5438 5430
rect 5846 5428 5880 5430
rect 6104 5428 6138 5430
rect 6546 5428 6580 5430
rect 6804 5428 6838 5430
rect 7246 5428 7280 5430
rect 7504 5428 7538 5430
rect 7946 5428 7980 5430
rect 8204 5428 8238 5430
rect 8646 5428 8680 5430
rect 8904 5428 8938 5430
rect 9346 5428 9380 5430
rect 9604 5428 9638 5430
rect 10046 5428 10080 5430
rect 10304 5428 10338 5430
rect -1196 5404 -1162 5406
rect -754 5404 -720 5406
rect -496 5404 -462 5406
rect -54 5404 -20 5406
rect 204 5404 238 5406
rect 646 5404 680 5406
rect 904 5404 938 5406
rect 1346 5404 1380 5406
rect 1604 5404 1638 5406
rect 2046 5404 2080 5406
rect 2304 5404 2338 5406
rect 3746 5404 3780 5406
rect 4004 5404 4038 5406
rect 4446 5404 4480 5406
rect 4704 5404 4738 5406
rect 5146 5404 5180 5406
rect 5404 5404 5438 5406
rect 5846 5404 5880 5406
rect 6104 5404 6138 5406
rect 6546 5404 6580 5406
rect 6804 5404 6838 5406
rect 7246 5404 7280 5406
rect 7504 5404 7538 5406
rect 7946 5404 7980 5406
rect 8204 5404 8238 5406
rect 8646 5404 8680 5406
rect 8904 5404 8938 5406
rect 9346 5404 9380 5406
rect 9604 5404 9638 5406
rect 10046 5404 10080 5406
rect 10304 5404 10338 5406
rect 11832 5405 12038 5539
rect 12732 5405 12938 5539
rect 13632 5405 13838 5539
rect 14532 5405 14738 5539
rect 15432 5405 15587 5539
rect -1196 5366 -1162 5368
rect -754 5366 -720 5368
rect -496 5366 -462 5368
rect -54 5366 -20 5368
rect 204 5366 238 5368
rect 646 5366 680 5368
rect 904 5366 938 5368
rect 1346 5366 1380 5368
rect 1604 5366 1638 5368
rect 2046 5366 2080 5368
rect 2304 5366 2338 5368
rect 3746 5366 3780 5368
rect 4004 5366 4038 5368
rect 4446 5366 4480 5368
rect 4704 5366 4738 5368
rect 5146 5366 5180 5368
rect 5404 5366 5438 5368
rect 5846 5366 5880 5368
rect 6104 5366 6138 5368
rect 6546 5366 6580 5368
rect 6804 5366 6838 5368
rect 7246 5366 7280 5368
rect 7504 5366 7538 5368
rect 7946 5366 7980 5368
rect 8204 5366 8238 5368
rect 8646 5366 8680 5368
rect 8904 5366 8938 5368
rect 9346 5366 9380 5368
rect 9604 5366 9638 5368
rect 10046 5366 10080 5368
rect 10304 5366 10338 5368
rect -1196 5360 -1162 5362
rect -754 5360 -720 5362
rect -496 5360 -462 5362
rect -54 5360 -20 5362
rect 204 5360 238 5362
rect 646 5360 680 5362
rect 904 5360 938 5362
rect 1346 5360 1380 5362
rect 1604 5360 1638 5362
rect 2046 5360 2080 5362
rect 2304 5360 2338 5362
rect 3746 5360 3780 5362
rect 4004 5360 4038 5362
rect 4446 5360 4480 5362
rect 4704 5360 4738 5362
rect 5146 5360 5180 5362
rect 5404 5360 5438 5362
rect 5846 5360 5880 5362
rect 6104 5360 6138 5362
rect 6546 5360 6580 5362
rect 6804 5360 6838 5362
rect 7246 5360 7280 5362
rect 7504 5360 7538 5362
rect 7946 5360 7980 5362
rect 8204 5360 8238 5362
rect 8646 5360 8680 5362
rect 8904 5360 8938 5362
rect 9346 5360 9380 5362
rect 9604 5360 9638 5362
rect 10046 5360 10080 5362
rect 10304 5360 10338 5362
rect -1196 5332 -1162 5334
rect -754 5332 -720 5334
rect -496 5332 -462 5334
rect -54 5332 -20 5334
rect 204 5332 238 5334
rect 646 5332 680 5334
rect 904 5332 938 5334
rect 1346 5332 1380 5334
rect 1604 5332 1638 5334
rect 2046 5332 2080 5334
rect 2304 5332 2338 5334
rect 3746 5332 3780 5334
rect 4004 5332 4038 5334
rect 4446 5332 4480 5334
rect 4704 5332 4738 5334
rect 5146 5332 5180 5334
rect 5404 5332 5438 5334
rect 5846 5332 5880 5334
rect 6104 5332 6138 5334
rect 6546 5332 6580 5334
rect 6804 5332 6838 5334
rect 7246 5332 7280 5334
rect 7504 5332 7538 5334
rect 7946 5332 7980 5334
rect 8204 5332 8238 5334
rect 8646 5332 8680 5334
rect 8904 5332 8938 5334
rect 9346 5332 9380 5334
rect 9604 5332 9638 5334
rect 10046 5332 10080 5334
rect 10304 5332 10338 5334
rect -1196 5292 -1162 5296
rect -754 5292 -720 5296
rect -496 5292 -462 5296
rect -54 5292 -20 5296
rect 204 5292 238 5296
rect 646 5292 680 5296
rect 904 5292 938 5296
rect 1346 5292 1380 5296
rect 1604 5292 1638 5296
rect 2046 5292 2080 5296
rect 2304 5292 2338 5296
rect 3746 5292 3780 5296
rect 4004 5292 4038 5296
rect 4446 5292 4480 5296
rect 4704 5292 4738 5296
rect 5146 5292 5180 5296
rect 5404 5292 5438 5296
rect 5846 5292 5880 5296
rect 6104 5292 6138 5296
rect 6546 5292 6580 5296
rect 6804 5292 6838 5296
rect 7246 5292 7280 5296
rect 7504 5292 7538 5296
rect 7946 5292 7980 5296
rect 8204 5292 8238 5296
rect 8646 5292 8680 5296
rect 8904 5292 8938 5296
rect 9346 5292 9380 5296
rect 9604 5292 9638 5296
rect 10046 5292 10080 5296
rect 10304 5292 10338 5296
rect -1196 5260 -1162 5262
rect -754 5260 -720 5262
rect -496 5260 -462 5262
rect -54 5260 -20 5262
rect 204 5260 238 5262
rect 646 5260 680 5262
rect 904 5260 938 5262
rect 1346 5260 1380 5262
rect 1604 5260 1638 5262
rect 2046 5260 2080 5262
rect 2304 5260 2338 5262
rect 3746 5260 3780 5262
rect 4004 5260 4038 5262
rect 4446 5260 4480 5262
rect 4704 5260 4738 5262
rect 5146 5260 5180 5262
rect 5404 5260 5438 5262
rect 5846 5260 5880 5262
rect 6104 5260 6138 5262
rect 6546 5260 6580 5262
rect 6804 5260 6838 5262
rect 7246 5260 7280 5262
rect 7504 5260 7538 5262
rect 7946 5260 7980 5262
rect 8204 5260 8238 5262
rect 8646 5260 8680 5262
rect 8904 5260 8938 5262
rect 9346 5260 9380 5262
rect 9604 5260 9638 5262
rect 10046 5260 10080 5262
rect 10304 5260 10338 5262
rect -1196 5222 -1162 5226
rect -754 5222 -720 5226
rect -496 5222 -462 5226
rect -54 5222 -20 5226
rect 204 5222 238 5226
rect 646 5222 680 5226
rect 904 5222 938 5226
rect 1346 5222 1380 5226
rect 1604 5222 1638 5226
rect 2046 5222 2080 5226
rect 2304 5222 2338 5226
rect 3746 5222 3780 5226
rect 4004 5222 4038 5226
rect 4446 5222 4480 5226
rect 4704 5222 4738 5226
rect 5146 5222 5180 5226
rect 5404 5222 5438 5226
rect 5846 5222 5880 5226
rect 6104 5222 6138 5226
rect 6546 5222 6580 5226
rect 6804 5222 6838 5226
rect 7246 5222 7280 5226
rect 7504 5222 7538 5226
rect 7946 5222 7980 5226
rect 8204 5222 8238 5226
rect 8646 5222 8680 5226
rect 8904 5222 8938 5226
rect 9346 5222 9380 5226
rect 9604 5222 9638 5226
rect 10046 5222 10080 5226
rect 10304 5222 10338 5226
rect -1196 5188 -1162 5190
rect -754 5188 -720 5190
rect -496 5188 -462 5190
rect -54 5188 -20 5190
rect 204 5188 238 5190
rect 646 5188 680 5190
rect 904 5188 938 5190
rect 1346 5188 1380 5190
rect 1604 5188 1638 5190
rect 2046 5188 2080 5190
rect 2304 5188 2338 5190
rect 3746 5188 3780 5190
rect 4004 5188 4038 5190
rect 4446 5188 4480 5190
rect 4704 5188 4738 5190
rect 5146 5188 5180 5190
rect 5404 5188 5438 5190
rect 5846 5188 5880 5190
rect 6104 5188 6138 5190
rect 6546 5188 6580 5190
rect 6804 5188 6838 5190
rect 7246 5188 7280 5190
rect 7504 5188 7538 5190
rect 7946 5188 7980 5190
rect 8204 5188 8238 5190
rect 8646 5188 8680 5190
rect 8904 5188 8938 5190
rect 9346 5188 9380 5190
rect 9604 5188 9638 5190
rect 10046 5188 10080 5190
rect 10304 5188 10338 5190
rect -1196 5156 -1162 5158
rect -754 5156 -720 5158
rect -496 5156 -462 5158
rect -54 5156 -20 5158
rect 204 5156 238 5158
rect 646 5156 680 5158
rect 904 5156 938 5158
rect 1346 5156 1380 5158
rect 1604 5156 1638 5158
rect 2046 5156 2080 5158
rect 2304 5156 2338 5158
rect 3746 5156 3780 5158
rect 4004 5156 4038 5158
rect 4446 5156 4480 5158
rect 4704 5156 4738 5158
rect 5146 5156 5180 5158
rect 5404 5156 5438 5158
rect 5846 5156 5880 5158
rect 6104 5156 6138 5158
rect 6546 5156 6580 5158
rect 6804 5156 6838 5158
rect 7246 5156 7280 5158
rect 7504 5156 7538 5158
rect 7946 5156 7980 5158
rect 8204 5156 8238 5158
rect 8646 5156 8680 5158
rect 8904 5156 8938 5158
rect 9346 5156 9380 5158
rect 9604 5156 9638 5158
rect 10046 5156 10080 5158
rect 10304 5156 10338 5158
rect -1196 5150 -1162 5152
rect -754 5150 -720 5152
rect -496 5150 -462 5152
rect -54 5150 -20 5152
rect 204 5150 238 5152
rect 646 5150 680 5152
rect 904 5150 938 5152
rect 1346 5150 1380 5152
rect 1604 5150 1638 5152
rect 2046 5150 2080 5152
rect 2304 5150 2338 5152
rect 3746 5150 3780 5152
rect 4004 5150 4038 5152
rect 4446 5150 4480 5152
rect 4704 5150 4738 5152
rect 5146 5150 5180 5152
rect 5404 5150 5438 5152
rect 5846 5150 5880 5152
rect 6104 5150 6138 5152
rect 6546 5150 6580 5152
rect 6804 5150 6838 5152
rect 7246 5150 7280 5152
rect 7504 5150 7538 5152
rect 7946 5150 7980 5152
rect 8204 5150 8238 5152
rect 8646 5150 8680 5152
rect 8904 5150 8938 5152
rect 9346 5150 9380 5152
rect 9604 5150 9638 5152
rect 10046 5150 10080 5152
rect 10304 5150 10338 5152
rect -1196 5116 -1162 5118
rect -754 5116 -720 5118
rect -496 5116 -462 5118
rect -54 5116 -20 5118
rect 204 5116 238 5118
rect 646 5116 680 5118
rect 904 5116 938 5118
rect 1346 5116 1380 5118
rect 1604 5116 1638 5118
rect 2046 5116 2080 5118
rect 2304 5116 2338 5118
rect 3746 5116 3780 5118
rect 4004 5116 4038 5118
rect 4446 5116 4480 5118
rect 4704 5116 4738 5118
rect 5146 5116 5180 5118
rect 5404 5116 5438 5118
rect 5846 5116 5880 5118
rect 6104 5116 6138 5118
rect 6546 5116 6580 5118
rect 6804 5116 6838 5118
rect 7246 5116 7280 5118
rect 7504 5116 7538 5118
rect 7946 5116 7980 5118
rect 8204 5116 8238 5118
rect 8646 5116 8680 5118
rect 8904 5116 8938 5118
rect 9346 5116 9380 5118
rect 9604 5116 9638 5118
rect 10046 5116 10080 5118
rect 10304 5116 10338 5118
rect -1196 5088 -1162 5090
rect -754 5088 -720 5090
rect -496 5088 -462 5090
rect -54 5088 -20 5090
rect 204 5088 238 5090
rect 646 5088 680 5090
rect 904 5088 938 5090
rect 1346 5088 1380 5090
rect 1604 5088 1638 5090
rect 2046 5088 2080 5090
rect 2304 5088 2338 5090
rect 3746 5088 3780 5090
rect 4004 5088 4038 5090
rect 4446 5088 4480 5090
rect 4704 5088 4738 5090
rect 5146 5088 5180 5090
rect 5404 5088 5438 5090
rect 5846 5088 5880 5090
rect 6104 5088 6138 5090
rect 6546 5088 6580 5090
rect 6804 5088 6838 5090
rect 7246 5088 7280 5090
rect 7504 5088 7538 5090
rect 7946 5088 7980 5090
rect 8204 5088 8238 5090
rect 8646 5088 8680 5090
rect 8904 5088 8938 5090
rect 9346 5088 9380 5090
rect 9604 5088 9638 5090
rect 10046 5088 10080 5090
rect 10304 5088 10338 5090
rect -1196 5078 -1162 5080
rect -754 5078 -720 5080
rect -496 5078 -462 5080
rect -54 5078 -20 5080
rect 204 5078 238 5080
rect 646 5078 680 5080
rect 904 5078 938 5080
rect 1346 5078 1380 5080
rect 1604 5078 1638 5080
rect 2046 5078 2080 5080
rect 2304 5078 2338 5080
rect 3746 5078 3780 5080
rect 4004 5078 4038 5080
rect 4446 5078 4480 5080
rect 4704 5078 4738 5080
rect 5146 5078 5180 5080
rect 5404 5078 5438 5080
rect 5846 5078 5880 5080
rect 6104 5078 6138 5080
rect 6546 5078 6580 5080
rect 6804 5078 6838 5080
rect 7246 5078 7280 5080
rect 7504 5078 7538 5080
rect 7946 5078 7980 5080
rect 8204 5078 8238 5080
rect 8646 5078 8680 5080
rect 8904 5078 8938 5080
rect 9346 5078 9380 5080
rect 9604 5078 9638 5080
rect 10046 5078 10080 5080
rect 10304 5078 10338 5080
rect -1196 5044 -1162 5046
rect -754 5044 -720 5046
rect -496 5044 -462 5046
rect -54 5044 -20 5046
rect 204 5044 238 5046
rect 646 5044 680 5046
rect 904 5044 938 5046
rect 1346 5044 1380 5046
rect 1604 5044 1638 5046
rect 2046 5044 2080 5046
rect 2304 5044 2338 5046
rect 3746 5044 3780 5046
rect 4004 5044 4038 5046
rect 4446 5044 4480 5046
rect 4704 5044 4738 5046
rect 5146 5044 5180 5046
rect 5404 5044 5438 5046
rect 5846 5044 5880 5046
rect 6104 5044 6138 5046
rect 6546 5044 6580 5046
rect 6804 5044 6838 5046
rect 7246 5044 7280 5046
rect 7504 5044 7538 5046
rect 7946 5044 7980 5046
rect 8204 5044 8238 5046
rect 8646 5044 8680 5046
rect 8904 5044 8938 5046
rect 9346 5044 9380 5046
rect 9604 5044 9638 5046
rect 10046 5044 10080 5046
rect 10304 5044 10338 5046
rect -1196 5020 -1162 5022
rect -754 5020 -720 5022
rect -496 5020 -462 5022
rect -54 5020 -20 5022
rect 204 5020 238 5022
rect 646 5020 680 5022
rect 904 5020 938 5022
rect 1346 5020 1380 5022
rect 1604 5020 1638 5022
rect 2046 5020 2080 5022
rect 2304 5020 2338 5022
rect 3746 5020 3780 5022
rect 4004 5020 4038 5022
rect 4446 5020 4480 5022
rect 4704 5020 4738 5022
rect 5146 5020 5180 5022
rect 5404 5020 5438 5022
rect 5846 5020 5880 5022
rect 6104 5020 6138 5022
rect 6546 5020 6580 5022
rect 6804 5020 6838 5022
rect 7246 5020 7280 5022
rect 7504 5020 7538 5022
rect 7946 5020 7980 5022
rect 8204 5020 8238 5022
rect 8646 5020 8680 5022
rect 8904 5020 8938 5022
rect 9346 5020 9380 5022
rect 9604 5020 9638 5022
rect 10046 5020 10080 5022
rect 10304 5020 10338 5022
rect -1196 5006 -1162 5008
rect -754 5006 -720 5008
rect -496 5006 -462 5008
rect -54 5006 -20 5008
rect 204 5006 238 5008
rect 646 5006 680 5008
rect 904 5006 938 5008
rect 1346 5006 1380 5008
rect 1604 5006 1638 5008
rect 2046 5006 2080 5008
rect 2304 5006 2338 5008
rect 3746 5006 3780 5008
rect 4004 5006 4038 5008
rect 4446 5006 4480 5008
rect 4704 5006 4738 5008
rect 5146 5006 5180 5008
rect 5404 5006 5438 5008
rect 5846 5006 5880 5008
rect 6104 5006 6138 5008
rect 6546 5006 6580 5008
rect 6804 5006 6838 5008
rect 7246 5006 7280 5008
rect 7504 5006 7538 5008
rect 7946 5006 7980 5008
rect 8204 5006 8238 5008
rect 8646 5006 8680 5008
rect 8904 5006 8938 5008
rect 9346 5006 9380 5008
rect 9604 5006 9638 5008
rect 10046 5006 10080 5008
rect 10304 5006 10338 5008
rect -1196 4972 -1162 4974
rect -754 4972 -720 4974
rect -496 4972 -462 4974
rect -54 4972 -20 4974
rect 204 4972 238 4974
rect 646 4972 680 4974
rect 904 4972 938 4974
rect 1346 4972 1380 4974
rect 1604 4972 1638 4974
rect 2046 4972 2080 4974
rect 2304 4972 2338 4974
rect 3746 4972 3780 4974
rect 4004 4972 4038 4974
rect 4446 4972 4480 4974
rect 4704 4972 4738 4974
rect 5146 4972 5180 4974
rect 5404 4972 5438 4974
rect 5846 4972 5880 4974
rect 6104 4972 6138 4974
rect 6546 4972 6580 4974
rect 6804 4972 6838 4974
rect 7246 4972 7280 4974
rect 7504 4972 7538 4974
rect 7946 4972 7980 4974
rect 8204 4972 8238 4974
rect 8646 4972 8680 4974
rect 8904 4972 8938 4974
rect 9346 4972 9380 4974
rect 9604 4972 9638 4974
rect 10046 4972 10080 4974
rect 10304 4972 10338 4974
rect -1196 4952 -1162 4954
rect -754 4952 -720 4954
rect -496 4952 -462 4954
rect -54 4952 -20 4954
rect 204 4952 238 4954
rect 646 4952 680 4954
rect 904 4952 938 4954
rect 1346 4952 1380 4954
rect 1604 4952 1638 4954
rect 2046 4952 2080 4954
rect 2304 4952 2338 4954
rect 3746 4952 3780 4954
rect 4004 4952 4038 4954
rect 4446 4952 4480 4954
rect 4704 4952 4738 4954
rect 5146 4952 5180 4954
rect 5404 4952 5438 4954
rect 5846 4952 5880 4954
rect 6104 4952 6138 4954
rect 6546 4952 6580 4954
rect 6804 4952 6838 4954
rect 7246 4952 7280 4954
rect 7504 4952 7538 4954
rect 7946 4952 7980 4954
rect 8204 4952 8238 4954
rect 8646 4952 8680 4954
rect 8904 4952 8938 4954
rect 9346 4952 9380 4954
rect 9604 4952 9638 4954
rect 10046 4952 10080 4954
rect 10304 4952 10338 4954
rect -1196 4934 -1162 4936
rect -754 4934 -720 4936
rect -496 4934 -462 4936
rect -54 4934 -20 4936
rect 204 4934 238 4936
rect 646 4934 680 4936
rect 904 4934 938 4936
rect 1346 4934 1380 4936
rect 1604 4934 1638 4936
rect 2046 4934 2080 4936
rect 2304 4934 2338 4936
rect 3746 4934 3780 4936
rect 4004 4934 4038 4936
rect 4446 4934 4480 4936
rect 4704 4934 4738 4936
rect 5146 4934 5180 4936
rect 5404 4934 5438 4936
rect 5846 4934 5880 4936
rect 6104 4934 6138 4936
rect 6546 4934 6580 4936
rect 6804 4934 6838 4936
rect 7246 4934 7280 4936
rect 7504 4934 7538 4936
rect 7946 4934 7980 4936
rect 8204 4934 8238 4936
rect 8646 4934 8680 4936
rect 8904 4934 8938 4936
rect 9346 4934 9380 4936
rect 9604 4934 9638 4936
rect 10046 4934 10080 4936
rect 10304 4934 10338 4936
rect -1196 4900 -1162 4902
rect -754 4900 -720 4902
rect -496 4900 -462 4902
rect -54 4900 -20 4902
rect 204 4900 238 4902
rect 646 4900 680 4902
rect 904 4900 938 4902
rect 1346 4900 1380 4902
rect 1604 4900 1638 4902
rect 2046 4900 2080 4902
rect 2304 4900 2338 4902
rect 3746 4900 3780 4902
rect 4004 4900 4038 4902
rect 4446 4900 4480 4902
rect 4704 4900 4738 4902
rect 5146 4900 5180 4902
rect 5404 4900 5438 4902
rect 5846 4900 5880 4902
rect 6104 4900 6138 4902
rect 6546 4900 6580 4902
rect 6804 4900 6838 4902
rect 7246 4900 7280 4902
rect 7504 4900 7538 4902
rect 7946 4900 7980 4902
rect 8204 4900 8238 4902
rect 8646 4900 8680 4902
rect 8904 4900 8938 4902
rect 9346 4900 9380 4902
rect 9604 4900 9638 4902
rect 10046 4900 10080 4902
rect 10304 4900 10338 4902
rect -1196 4884 -1162 4886
rect -754 4884 -720 4886
rect -496 4884 -462 4886
rect -54 4884 -20 4886
rect 204 4884 238 4886
rect 646 4884 680 4886
rect 904 4884 938 4886
rect 1346 4884 1380 4886
rect 1604 4884 1638 4886
rect 2046 4884 2080 4886
rect 2304 4884 2338 4886
rect 3746 4884 3780 4886
rect 4004 4884 4038 4886
rect 4446 4884 4480 4886
rect 4704 4884 4738 4886
rect 5146 4884 5180 4886
rect 5404 4884 5438 4886
rect 5846 4884 5880 4886
rect 6104 4884 6138 4886
rect 6546 4884 6580 4886
rect 6804 4884 6838 4886
rect 7246 4884 7280 4886
rect 7504 4884 7538 4886
rect 7946 4884 7980 4886
rect 8204 4884 8238 4886
rect 8646 4884 8680 4886
rect 8904 4884 8938 4886
rect 9346 4884 9380 4886
rect 9604 4884 9638 4886
rect 10046 4884 10080 4886
rect 10304 4884 10338 4886
rect -1196 4862 -1162 4864
rect -754 4862 -720 4864
rect -496 4862 -462 4864
rect -54 4862 -20 4864
rect 204 4862 238 4864
rect 646 4862 680 4864
rect 904 4862 938 4864
rect 1346 4862 1380 4864
rect 1604 4862 1638 4864
rect 2046 4862 2080 4864
rect 2304 4862 2338 4864
rect 3746 4862 3780 4864
rect 4004 4862 4038 4864
rect 4446 4862 4480 4864
rect 4704 4862 4738 4864
rect 5146 4862 5180 4864
rect 5404 4862 5438 4864
rect 5846 4862 5880 4864
rect 6104 4862 6138 4864
rect 6546 4862 6580 4864
rect 6804 4862 6838 4864
rect 7246 4862 7280 4864
rect 7504 4862 7538 4864
rect 7946 4862 7980 4864
rect 8204 4862 8238 4864
rect 8646 4862 8680 4864
rect 8904 4862 8938 4864
rect 9346 4862 9380 4864
rect 9604 4862 9638 4864
rect 10046 4862 10080 4864
rect 10304 4862 10338 4864
rect -1196 4828 -1162 4830
rect -754 4828 -720 4830
rect -496 4828 -462 4830
rect -54 4828 -20 4830
rect 204 4828 238 4830
rect 646 4828 680 4830
rect 904 4828 938 4830
rect 1346 4828 1380 4830
rect 1604 4828 1638 4830
rect 2046 4828 2080 4830
rect 2304 4828 2338 4830
rect 3746 4828 3780 4830
rect 4004 4828 4038 4830
rect 4446 4828 4480 4830
rect 4704 4828 4738 4830
rect 5146 4828 5180 4830
rect 5404 4828 5438 4830
rect 5846 4828 5880 4830
rect 6104 4828 6138 4830
rect 6546 4828 6580 4830
rect 6804 4828 6838 4830
rect 7246 4828 7280 4830
rect 7504 4828 7538 4830
rect 7946 4828 7980 4830
rect 8204 4828 8238 4830
rect 8646 4828 8680 4830
rect 8904 4828 8938 4830
rect 9346 4828 9380 4830
rect 9604 4828 9638 4830
rect 10046 4828 10080 4830
rect 10304 4828 10338 4830
rect -1196 4816 -1162 4818
rect -754 4816 -720 4818
rect -496 4816 -462 4818
rect -54 4816 -20 4818
rect 204 4816 238 4818
rect 646 4816 680 4818
rect 904 4816 938 4818
rect 1346 4816 1380 4818
rect 1604 4816 1638 4818
rect 2046 4816 2080 4818
rect 2304 4816 2338 4818
rect 3746 4816 3780 4818
rect 4004 4816 4038 4818
rect 4446 4816 4480 4818
rect 4704 4816 4738 4818
rect 5146 4816 5180 4818
rect 5404 4816 5438 4818
rect 5846 4816 5880 4818
rect 6104 4816 6138 4818
rect 6546 4816 6580 4818
rect 6804 4816 6838 4818
rect 7246 4816 7280 4818
rect 7504 4816 7538 4818
rect 7946 4816 7980 4818
rect 8204 4816 8238 4818
rect 8646 4816 8680 4818
rect 8904 4816 8938 4818
rect 9346 4816 9380 4818
rect 9604 4816 9638 4818
rect 10046 4816 10080 4818
rect 10304 4816 10338 4818
rect -1196 4790 -1162 4792
rect -754 4790 -720 4792
rect -496 4790 -462 4792
rect -54 4790 -20 4792
rect 204 4790 238 4792
rect 646 4790 680 4792
rect 904 4790 938 4792
rect 1346 4790 1380 4792
rect 1604 4790 1638 4792
rect 2046 4790 2080 4792
rect 2304 4790 2338 4792
rect 3746 4790 3780 4792
rect 4004 4790 4038 4792
rect 4446 4790 4480 4792
rect 4704 4790 4738 4792
rect 5146 4790 5180 4792
rect 5404 4790 5438 4792
rect 5846 4790 5880 4792
rect 6104 4790 6138 4792
rect 6546 4790 6580 4792
rect 6804 4790 6838 4792
rect 7246 4790 7280 4792
rect 7504 4790 7538 4792
rect 7946 4790 7980 4792
rect 8204 4790 8238 4792
rect 8646 4790 8680 4792
rect 8904 4790 8938 4792
rect 9346 4790 9380 4792
rect 9604 4790 9638 4792
rect 10046 4790 10080 4792
rect 10304 4790 10338 4792
rect -1196 4756 -1162 4758
rect -754 4756 -720 4758
rect -496 4756 -462 4758
rect -54 4756 -20 4758
rect 204 4756 238 4758
rect 646 4756 680 4758
rect 904 4756 938 4758
rect 1346 4756 1380 4758
rect 1604 4756 1638 4758
rect 2046 4756 2080 4758
rect 2304 4756 2338 4758
rect 3746 4756 3780 4758
rect 4004 4756 4038 4758
rect 4446 4756 4480 4758
rect 4704 4756 4738 4758
rect 5146 4756 5180 4758
rect 5404 4756 5438 4758
rect 5846 4756 5880 4758
rect 6104 4756 6138 4758
rect 6546 4756 6580 4758
rect 6804 4756 6838 4758
rect 7246 4756 7280 4758
rect 7504 4756 7538 4758
rect 7946 4756 7980 4758
rect 8204 4756 8238 4758
rect 8646 4756 8680 4758
rect 8904 4756 8938 4758
rect 9346 4756 9380 4758
rect 9604 4756 9638 4758
rect 10046 4756 10080 4758
rect 10304 4756 10338 4758
rect -1196 4748 -1162 4750
rect -754 4748 -720 4750
rect -496 4748 -462 4750
rect -54 4748 -20 4750
rect 204 4748 238 4750
rect 646 4748 680 4750
rect 904 4748 938 4750
rect 1346 4748 1380 4750
rect 1604 4748 1638 4750
rect 2046 4748 2080 4750
rect 2304 4748 2338 4750
rect 3746 4748 3780 4750
rect 4004 4748 4038 4750
rect 4446 4748 4480 4750
rect 4704 4748 4738 4750
rect 5146 4748 5180 4750
rect 5404 4748 5438 4750
rect 5846 4748 5880 4750
rect 6104 4748 6138 4750
rect 6546 4748 6580 4750
rect 6804 4748 6838 4750
rect 7246 4748 7280 4750
rect 7504 4748 7538 4750
rect 7946 4748 7980 4750
rect 8204 4748 8238 4750
rect 8646 4748 8680 4750
rect 8904 4748 8938 4750
rect 9346 4748 9380 4750
rect 9604 4748 9638 4750
rect 10046 4748 10080 4750
rect 10304 4748 10338 4750
rect -1196 4718 -1162 4720
rect -754 4718 -720 4720
rect -496 4718 -462 4720
rect -54 4718 -20 4720
rect 204 4718 238 4720
rect 646 4718 680 4720
rect 904 4718 938 4720
rect 1346 4718 1380 4720
rect 1604 4718 1638 4720
rect 2046 4718 2080 4720
rect 2304 4718 2338 4720
rect 3746 4718 3780 4720
rect 4004 4718 4038 4720
rect 4446 4718 4480 4720
rect 4704 4718 4738 4720
rect 5146 4718 5180 4720
rect 5404 4718 5438 4720
rect 5846 4718 5880 4720
rect 6104 4718 6138 4720
rect 6546 4718 6580 4720
rect 6804 4718 6838 4720
rect 7246 4718 7280 4720
rect 7504 4718 7538 4720
rect 7946 4718 7980 4720
rect 8204 4718 8238 4720
rect 8646 4718 8680 4720
rect 8904 4718 8938 4720
rect 9346 4718 9380 4720
rect 9604 4718 9638 4720
rect 10046 4718 10080 4720
rect 10304 4718 10338 4720
rect -1196 4684 -1162 4686
rect -754 4684 -720 4686
rect -496 4684 -462 4686
rect -54 4684 -20 4686
rect 204 4684 238 4686
rect 646 4684 680 4686
rect 904 4684 938 4686
rect 1346 4684 1380 4686
rect 1604 4684 1638 4686
rect 2046 4684 2080 4686
rect 2304 4684 2338 4686
rect 3746 4684 3780 4686
rect 4004 4684 4038 4686
rect 4446 4684 4480 4686
rect 4704 4684 4738 4686
rect 5146 4684 5180 4686
rect 5404 4684 5438 4686
rect 5846 4684 5880 4686
rect 6104 4684 6138 4686
rect 6546 4684 6580 4686
rect 6804 4684 6838 4686
rect 7246 4684 7280 4686
rect 7504 4684 7538 4686
rect 7946 4684 7980 4686
rect 8204 4684 8238 4686
rect 8646 4684 8680 4686
rect 8904 4684 8938 4686
rect 9346 4684 9380 4686
rect 9604 4684 9638 4686
rect 10046 4684 10080 4686
rect 10304 4684 10338 4686
rect -1196 4680 -1162 4682
rect -754 4680 -720 4682
rect -496 4680 -462 4682
rect -54 4680 -20 4682
rect 204 4680 238 4682
rect 646 4680 680 4682
rect 904 4680 938 4682
rect 1346 4680 1380 4682
rect 1604 4680 1638 4682
rect 2046 4680 2080 4682
rect 2304 4680 2338 4682
rect 3746 4680 3780 4682
rect 4004 4680 4038 4682
rect 4446 4680 4480 4682
rect 4704 4680 4738 4682
rect 5146 4680 5180 4682
rect 5404 4680 5438 4682
rect 5846 4680 5880 4682
rect 6104 4680 6138 4682
rect 6546 4680 6580 4682
rect 6804 4680 6838 4682
rect 7246 4680 7280 4682
rect 7504 4680 7538 4682
rect 7946 4680 7980 4682
rect 8204 4680 8238 4682
rect 8646 4680 8680 4682
rect 8904 4680 8938 4682
rect 9346 4680 9380 4682
rect 9604 4680 9638 4682
rect 10046 4680 10080 4682
rect 10304 4680 10338 4682
rect -1196 4646 -1162 4648
rect -754 4646 -720 4648
rect -496 4646 -462 4648
rect -54 4646 -20 4648
rect 204 4646 238 4648
rect 646 4646 680 4648
rect 904 4646 938 4648
rect 1346 4646 1380 4648
rect 1604 4646 1638 4648
rect 2046 4646 2080 4648
rect 2304 4646 2338 4648
rect 3746 4646 3780 4648
rect 4004 4646 4038 4648
rect 4446 4646 4480 4648
rect 4704 4646 4738 4648
rect 5146 4646 5180 4648
rect 5404 4646 5438 4648
rect 5846 4646 5880 4648
rect 6104 4646 6138 4648
rect 6546 4646 6580 4648
rect 6804 4646 6838 4648
rect 7246 4646 7280 4648
rect 7504 4646 7538 4648
rect 7946 4646 7980 4648
rect 8204 4646 8238 4648
rect 8646 4646 8680 4648
rect 8904 4646 8938 4648
rect 9346 4646 9380 4648
rect 9604 4646 9638 4648
rect 10046 4646 10080 4648
rect 10304 4646 10338 4648
rect -1196 4612 -1162 4614
rect -754 4612 -720 4614
rect -496 4612 -462 4614
rect -54 4612 -20 4614
rect 204 4612 238 4614
rect 646 4612 680 4614
rect 904 4612 938 4614
rect 1346 4612 1380 4614
rect 1604 4612 1638 4614
rect 2046 4612 2080 4614
rect 2304 4612 2338 4614
rect 3746 4612 3780 4614
rect 4004 4612 4038 4614
rect 4446 4612 4480 4614
rect 4704 4612 4738 4614
rect 5146 4612 5180 4614
rect 5404 4612 5438 4614
rect 5846 4612 5880 4614
rect 6104 4612 6138 4614
rect 6546 4612 6580 4614
rect 6804 4612 6838 4614
rect 7246 4612 7280 4614
rect 7504 4612 7538 4614
rect 7946 4612 7980 4614
rect 8204 4612 8238 4614
rect 8646 4612 8680 4614
rect 8904 4612 8938 4614
rect 9346 4612 9380 4614
rect 9604 4612 9638 4614
rect 10046 4612 10080 4614
rect 10304 4612 10338 4614
rect -1196 4574 -1162 4576
rect -754 4574 -720 4576
rect -496 4574 -462 4576
rect -54 4574 -20 4576
rect 204 4574 238 4576
rect 646 4574 680 4576
rect 904 4574 938 4576
rect 1346 4574 1380 4576
rect 1604 4574 1638 4576
rect 2046 4574 2080 4576
rect 2304 4574 2338 4576
rect 3746 4574 3780 4576
rect 4004 4574 4038 4576
rect 4446 4574 4480 4576
rect 4704 4574 4738 4576
rect 5146 4574 5180 4576
rect 5404 4574 5438 4576
rect 5846 4574 5880 4576
rect 6104 4574 6138 4576
rect 6546 4574 6580 4576
rect 6804 4574 6838 4576
rect 7246 4574 7280 4576
rect 7504 4574 7538 4576
rect 7946 4574 7980 4576
rect 8204 4574 8238 4576
rect 8646 4574 8680 4576
rect 8904 4574 8938 4576
rect 9346 4574 9380 4576
rect 9604 4574 9638 4576
rect 10046 4574 10080 4576
rect 10304 4574 10338 4576
rect -1196 4544 -1162 4546
rect -754 4544 -720 4546
rect -496 4544 -462 4546
rect -54 4544 -20 4546
rect 204 4544 238 4546
rect 646 4544 680 4546
rect 904 4544 938 4546
rect 1346 4544 1380 4546
rect 1604 4544 1638 4546
rect 2046 4544 2080 4546
rect 2304 4544 2338 4546
rect 3746 4544 3780 4546
rect 4004 4544 4038 4546
rect 4446 4544 4480 4546
rect 4704 4544 4738 4546
rect 5146 4544 5180 4546
rect 5404 4544 5438 4546
rect 5846 4544 5880 4546
rect 6104 4544 6138 4546
rect 6546 4544 6580 4546
rect 6804 4544 6838 4546
rect 7246 4544 7280 4546
rect 7504 4544 7538 4546
rect 7946 4544 7980 4546
rect 8204 4544 8238 4546
rect 8646 4544 8680 4546
rect 8904 4544 8938 4546
rect 9346 4544 9380 4546
rect 9604 4544 9638 4546
rect 10046 4544 10080 4546
rect 10304 4544 10338 4546
rect -1196 4540 -1162 4542
rect -754 4540 -720 4542
rect -496 4540 -462 4542
rect -54 4540 -20 4542
rect 204 4540 238 4542
rect 646 4540 680 4542
rect 904 4540 938 4542
rect 1346 4540 1380 4542
rect 1604 4540 1638 4542
rect 2046 4540 2080 4542
rect 2304 4540 2338 4542
rect 3746 4540 3780 4542
rect 4004 4540 4038 4542
rect 4446 4540 4480 4542
rect 4704 4540 4738 4542
rect 5146 4540 5180 4542
rect 5404 4540 5438 4542
rect 5846 4540 5880 4542
rect 6104 4540 6138 4542
rect 6546 4540 6580 4542
rect 6804 4540 6838 4542
rect 7246 4540 7280 4542
rect 7504 4540 7538 4542
rect 7946 4540 7980 4542
rect 8204 4540 8238 4542
rect 8646 4540 8680 4542
rect 8904 4540 8938 4542
rect 9346 4540 9380 4542
rect 9604 4540 9638 4542
rect 10046 4540 10080 4542
rect 10304 4540 10338 4542
rect -1196 4502 -1162 4504
rect -754 4502 -720 4504
rect -496 4502 -462 4504
rect -54 4502 -20 4504
rect 204 4502 238 4504
rect 646 4502 680 4504
rect 904 4502 938 4504
rect 1346 4502 1380 4504
rect 1604 4502 1638 4504
rect 2046 4502 2080 4504
rect 2304 4502 2338 4504
rect 3746 4502 3780 4504
rect 4004 4502 4038 4504
rect 4446 4502 4480 4504
rect 4704 4502 4738 4504
rect 5146 4502 5180 4504
rect 5404 4502 5438 4504
rect 5846 4502 5880 4504
rect 6104 4502 6138 4504
rect 6546 4502 6580 4504
rect 6804 4502 6838 4504
rect 7246 4502 7280 4504
rect 7504 4502 7538 4504
rect 7946 4502 7980 4504
rect 8204 4502 8238 4504
rect 8646 4502 8680 4504
rect 8904 4502 8938 4504
rect 9346 4502 9380 4504
rect 9604 4502 9638 4504
rect 10046 4502 10080 4504
rect 10304 4502 10338 4504
rect -1196 4476 -1162 4478
rect -754 4476 -720 4478
rect -496 4476 -462 4478
rect -54 4476 -20 4478
rect 204 4476 238 4478
rect 646 4476 680 4478
rect 904 4476 938 4478
rect 1346 4476 1380 4478
rect 1604 4476 1638 4478
rect 2046 4476 2080 4478
rect 2304 4476 2338 4478
rect 3746 4476 3780 4478
rect 4004 4476 4038 4478
rect 4446 4476 4480 4478
rect 4704 4476 4738 4478
rect 5146 4476 5180 4478
rect 5404 4476 5438 4478
rect 5846 4476 5880 4478
rect 6104 4476 6138 4478
rect 6546 4476 6580 4478
rect 6804 4476 6838 4478
rect 7246 4476 7280 4478
rect 7504 4476 7538 4478
rect 7946 4476 7980 4478
rect 8204 4476 8238 4478
rect 8646 4476 8680 4478
rect 8904 4476 8938 4478
rect 9346 4476 9380 4478
rect 9604 4476 9638 4478
rect 10046 4476 10080 4478
rect 10304 4476 10338 4478
rect -1196 4468 -1162 4470
rect -754 4468 -720 4470
rect -496 4468 -462 4470
rect -54 4468 -20 4470
rect 204 4468 238 4470
rect 646 4468 680 4470
rect 904 4468 938 4470
rect 1346 4468 1380 4470
rect 1604 4468 1638 4470
rect 2046 4468 2080 4470
rect 2304 4468 2338 4470
rect 3746 4468 3780 4470
rect 4004 4468 4038 4470
rect 4446 4468 4480 4470
rect 4704 4468 4738 4470
rect 5146 4468 5180 4470
rect 5404 4468 5438 4470
rect 5846 4468 5880 4470
rect 6104 4468 6138 4470
rect 6546 4468 6580 4470
rect 6804 4468 6838 4470
rect 7246 4468 7280 4470
rect 7504 4468 7538 4470
rect 7946 4468 7980 4470
rect 8204 4468 8238 4470
rect 8646 4468 8680 4470
rect 8904 4468 8938 4470
rect 9346 4468 9380 4470
rect 9604 4468 9638 4470
rect 10046 4468 10080 4470
rect 10304 4468 10338 4470
rect -1196 4430 -1162 4432
rect -754 4430 -720 4432
rect -496 4430 -462 4432
rect -54 4430 -20 4432
rect 204 4430 238 4432
rect 646 4430 680 4432
rect 904 4430 938 4432
rect 1346 4430 1380 4432
rect 1604 4430 1638 4432
rect 2046 4430 2080 4432
rect 2304 4430 2338 4432
rect 3746 4430 3780 4432
rect 4004 4430 4038 4432
rect 4446 4430 4480 4432
rect 4704 4430 4738 4432
rect 5146 4430 5180 4432
rect 5404 4430 5438 4432
rect 5846 4430 5880 4432
rect 6104 4430 6138 4432
rect 6546 4430 6580 4432
rect 6804 4430 6838 4432
rect 7246 4430 7280 4432
rect 7504 4430 7538 4432
rect 7946 4430 7980 4432
rect 8204 4430 8238 4432
rect 8646 4430 8680 4432
rect 8904 4430 8938 4432
rect 9346 4430 9380 4432
rect 9604 4430 9638 4432
rect 10046 4430 10080 4432
rect 10304 4430 10338 4432
rect -1196 4408 -1162 4410
rect -754 4408 -720 4410
rect -496 4408 -462 4410
rect -54 4408 -20 4410
rect 204 4408 238 4410
rect 646 4408 680 4410
rect 904 4408 938 4410
rect 1346 4408 1380 4410
rect 1604 4408 1638 4410
rect 2046 4408 2080 4410
rect 2304 4408 2338 4410
rect 3746 4408 3780 4410
rect 4004 4408 4038 4410
rect 4446 4408 4480 4410
rect 4704 4408 4738 4410
rect 5146 4408 5180 4410
rect 5404 4408 5438 4410
rect 5846 4408 5880 4410
rect 6104 4408 6138 4410
rect 6546 4408 6580 4410
rect 6804 4408 6838 4410
rect 7246 4408 7280 4410
rect 7504 4408 7538 4410
rect 7946 4408 7980 4410
rect 8204 4408 8238 4410
rect 8646 4408 8680 4410
rect 8904 4408 8938 4410
rect 9346 4408 9380 4410
rect 9604 4408 9638 4410
rect 10046 4408 10080 4410
rect 10304 4408 10338 4410
rect -1196 4396 -1162 4398
rect -754 4396 -720 4398
rect -496 4396 -462 4398
rect -54 4396 -20 4398
rect 204 4396 238 4398
rect 646 4396 680 4398
rect 904 4396 938 4398
rect 1346 4396 1380 4398
rect 1604 4396 1638 4398
rect 2046 4396 2080 4398
rect 2304 4396 2338 4398
rect 3746 4396 3780 4398
rect 4004 4396 4038 4398
rect 4446 4396 4480 4398
rect 4704 4396 4738 4398
rect 5146 4396 5180 4398
rect 5404 4396 5438 4398
rect 5846 4396 5880 4398
rect 6104 4396 6138 4398
rect 6546 4396 6580 4398
rect 6804 4396 6838 4398
rect 7246 4396 7280 4398
rect 7504 4396 7538 4398
rect 7946 4396 7980 4398
rect 8204 4396 8238 4398
rect 8646 4396 8680 4398
rect 8904 4396 8938 4398
rect 9346 4396 9380 4398
rect 9604 4396 9638 4398
rect 10046 4396 10080 4398
rect 10304 4396 10338 4398
rect -1196 4358 -1162 4360
rect -754 4358 -720 4360
rect -496 4358 -462 4360
rect -54 4358 -20 4360
rect 204 4358 238 4360
rect 646 4358 680 4360
rect 904 4358 938 4360
rect 1346 4358 1380 4360
rect 1604 4358 1638 4360
rect 2046 4358 2080 4360
rect 2304 4358 2338 4360
rect 3746 4358 3780 4360
rect 4004 4358 4038 4360
rect 4446 4358 4480 4360
rect 4704 4358 4738 4360
rect 5146 4358 5180 4360
rect 5404 4358 5438 4360
rect 5846 4358 5880 4360
rect 6104 4358 6138 4360
rect 6546 4358 6580 4360
rect 6804 4358 6838 4360
rect 7246 4358 7280 4360
rect 7504 4358 7538 4360
rect 7946 4358 7980 4360
rect 8204 4358 8238 4360
rect 8646 4358 8680 4360
rect 8904 4358 8938 4360
rect 9346 4358 9380 4360
rect 9604 4358 9638 4360
rect 10046 4358 10080 4360
rect 10304 4358 10338 4360
rect -1196 4340 -1162 4342
rect -754 4340 -720 4342
rect -496 4340 -462 4342
rect -54 4340 -20 4342
rect 204 4340 238 4342
rect 646 4340 680 4342
rect 904 4340 938 4342
rect 1346 4340 1380 4342
rect 1604 4340 1638 4342
rect 2046 4340 2080 4342
rect 2304 4340 2338 4342
rect 3746 4340 3780 4342
rect 4004 4340 4038 4342
rect 4446 4340 4480 4342
rect 4704 4340 4738 4342
rect 5146 4340 5180 4342
rect 5404 4340 5438 4342
rect 5846 4340 5880 4342
rect 6104 4340 6138 4342
rect 6546 4340 6580 4342
rect 6804 4340 6838 4342
rect 7246 4340 7280 4342
rect 7504 4340 7538 4342
rect 7946 4340 7980 4342
rect 8204 4340 8238 4342
rect 8646 4340 8680 4342
rect 8904 4340 8938 4342
rect 9346 4340 9380 4342
rect 9604 4340 9638 4342
rect 10046 4340 10080 4342
rect 10304 4340 10338 4342
rect -1196 4324 -1162 4326
rect -754 4324 -720 4326
rect -496 4324 -462 4326
rect -54 4324 -20 4326
rect 204 4324 238 4326
rect 646 4324 680 4326
rect 904 4324 938 4326
rect 1346 4324 1380 4326
rect 1604 4324 1638 4326
rect 2046 4324 2080 4326
rect 2304 4324 2338 4326
rect 3746 4324 3780 4326
rect 4004 4324 4038 4326
rect 4446 4324 4480 4326
rect 4704 4324 4738 4326
rect 5146 4324 5180 4326
rect 5404 4324 5438 4326
rect 5846 4324 5880 4326
rect 6104 4324 6138 4326
rect 6546 4324 6580 4326
rect 6804 4324 6838 4326
rect 7246 4324 7280 4326
rect 7504 4324 7538 4326
rect 7946 4324 7980 4326
rect 8204 4324 8238 4326
rect 8646 4324 8680 4326
rect 8904 4324 8938 4326
rect 9346 4324 9380 4326
rect 9604 4324 9638 4326
rect 10046 4324 10080 4326
rect 10304 4324 10338 4326
rect -1196 4286 -1162 4288
rect -754 4286 -720 4288
rect -496 4286 -462 4288
rect -54 4286 -20 4288
rect 204 4286 238 4288
rect 646 4286 680 4288
rect 904 4286 938 4288
rect 1346 4286 1380 4288
rect 1604 4286 1638 4288
rect 2046 4286 2080 4288
rect 2304 4286 2338 4288
rect 3746 4286 3780 4288
rect 4004 4286 4038 4288
rect 4446 4286 4480 4288
rect 4704 4286 4738 4288
rect 5146 4286 5180 4288
rect 5404 4286 5438 4288
rect 5846 4286 5880 4288
rect 6104 4286 6138 4288
rect 6546 4286 6580 4288
rect 6804 4286 6838 4288
rect 7246 4286 7280 4288
rect 7504 4286 7538 4288
rect 7946 4286 7980 4288
rect 8204 4286 8238 4288
rect 8646 4286 8680 4288
rect 8904 4286 8938 4288
rect 9346 4286 9380 4288
rect 9604 4286 9638 4288
rect 10046 4286 10080 4288
rect 10304 4286 10338 4288
rect -1196 4272 -1162 4274
rect -754 4272 -720 4274
rect -496 4272 -462 4274
rect -54 4272 -20 4274
rect 204 4272 238 4274
rect 646 4272 680 4274
rect 904 4272 938 4274
rect 1346 4272 1380 4274
rect 1604 4272 1638 4274
rect 2046 4272 2080 4274
rect 2304 4272 2338 4274
rect 3746 4272 3780 4274
rect 4004 4272 4038 4274
rect 4446 4272 4480 4274
rect 4704 4272 4738 4274
rect 5146 4272 5180 4274
rect 5404 4272 5438 4274
rect 5846 4272 5880 4274
rect 6104 4272 6138 4274
rect 6546 4272 6580 4274
rect 6804 4272 6838 4274
rect 7246 4272 7280 4274
rect 7504 4272 7538 4274
rect 7946 4272 7980 4274
rect 8204 4272 8238 4274
rect 8646 4272 8680 4274
rect 8904 4272 8938 4274
rect 9346 4272 9380 4274
rect 9604 4272 9638 4274
rect 10046 4272 10080 4274
rect 10304 4272 10338 4274
rect -1196 4252 -1162 4254
rect -754 4252 -720 4254
rect -496 4252 -462 4254
rect -54 4252 -20 4254
rect 204 4252 238 4254
rect 646 4252 680 4254
rect 904 4252 938 4254
rect 1346 4252 1380 4254
rect 1604 4252 1638 4254
rect 2046 4252 2080 4254
rect 2304 4252 2338 4254
rect 3746 4252 3780 4254
rect 4004 4252 4038 4254
rect 4446 4252 4480 4254
rect 4704 4252 4738 4254
rect 5146 4252 5180 4254
rect 5404 4252 5438 4254
rect 5846 4252 5880 4254
rect 6104 4252 6138 4254
rect 6546 4252 6580 4254
rect 6804 4252 6838 4254
rect 7246 4252 7280 4254
rect 7504 4252 7538 4254
rect 7946 4252 7980 4254
rect 8204 4252 8238 4254
rect 8646 4252 8680 4254
rect 8904 4252 8938 4254
rect 9346 4252 9380 4254
rect 9604 4252 9638 4254
rect 10046 4252 10080 4254
rect 10304 4252 10338 4254
rect -1196 4214 -1162 4216
rect -754 4214 -720 4216
rect -496 4214 -462 4216
rect -54 4214 -20 4216
rect 204 4214 238 4216
rect 646 4214 680 4216
rect 904 4214 938 4216
rect 1346 4214 1380 4216
rect 1604 4214 1638 4216
rect 2046 4214 2080 4216
rect 2304 4214 2338 4216
rect 3746 4214 3780 4216
rect 4004 4214 4038 4216
rect 4446 4214 4480 4216
rect 4704 4214 4738 4216
rect 5146 4214 5180 4216
rect 5404 4214 5438 4216
rect 5846 4214 5880 4216
rect 6104 4214 6138 4216
rect 6546 4214 6580 4216
rect 6804 4214 6838 4216
rect 7246 4214 7280 4216
rect 7504 4214 7538 4216
rect 7946 4214 7980 4216
rect 8204 4214 8238 4216
rect 8646 4214 8680 4216
rect 8904 4214 8938 4216
rect 9346 4214 9380 4216
rect 9604 4214 9638 4216
rect 10046 4214 10080 4216
rect 10304 4214 10338 4216
rect -1196 4204 -1162 4206
rect -754 4204 -720 4206
rect -496 4204 -462 4206
rect -54 4204 -20 4206
rect 204 4204 238 4206
rect 646 4204 680 4206
rect 904 4204 938 4206
rect 1346 4204 1380 4206
rect 1604 4204 1638 4206
rect 2046 4204 2080 4206
rect 2304 4204 2338 4206
rect 3746 4204 3780 4206
rect 4004 4204 4038 4206
rect 4446 4204 4480 4206
rect 4704 4204 4738 4206
rect 5146 4204 5180 4206
rect 5404 4204 5438 4206
rect 5846 4204 5880 4206
rect 6104 4204 6138 4206
rect 6546 4204 6580 4206
rect 6804 4204 6838 4206
rect 7246 4204 7280 4206
rect 7504 4204 7538 4206
rect 7946 4204 7980 4206
rect 8204 4204 8238 4206
rect 8646 4204 8680 4206
rect 8904 4204 8938 4206
rect 9346 4204 9380 4206
rect 9604 4204 9638 4206
rect 10046 4204 10080 4206
rect 10304 4204 10338 4206
rect -1196 4180 -1162 4182
rect -754 4180 -720 4182
rect -496 4180 -462 4182
rect -54 4180 -20 4182
rect 204 4180 238 4182
rect 646 4180 680 4182
rect 904 4180 938 4182
rect 1346 4180 1380 4182
rect 1604 4180 1638 4182
rect 2046 4180 2080 4182
rect 2304 4180 2338 4182
rect 3746 4180 3780 4182
rect 4004 4180 4038 4182
rect 4446 4180 4480 4182
rect 4704 4180 4738 4182
rect 5146 4180 5180 4182
rect 5404 4180 5438 4182
rect 5846 4180 5880 4182
rect 6104 4180 6138 4182
rect 6546 4180 6580 4182
rect 6804 4180 6838 4182
rect 7246 4180 7280 4182
rect 7504 4180 7538 4182
rect 7946 4180 7980 4182
rect 8204 4180 8238 4182
rect 8646 4180 8680 4182
rect 8904 4180 8938 4182
rect 9346 4180 9380 4182
rect 9604 4180 9638 4182
rect 10046 4180 10080 4182
rect 10304 4180 10338 4182
rect -1196 4142 -1162 4144
rect -754 4142 -720 4144
rect -496 4142 -462 4144
rect -54 4142 -20 4144
rect 204 4142 238 4144
rect 646 4142 680 4144
rect 904 4142 938 4144
rect 1346 4142 1380 4144
rect 1604 4142 1638 4144
rect 2046 4142 2080 4144
rect 2304 4142 2338 4144
rect 3746 4142 3780 4144
rect 4004 4142 4038 4144
rect 4446 4142 4480 4144
rect 4704 4142 4738 4144
rect 5146 4142 5180 4144
rect 5404 4142 5438 4144
rect 5846 4142 5880 4144
rect 6104 4142 6138 4144
rect 6546 4142 6580 4144
rect 6804 4142 6838 4144
rect 7246 4142 7280 4144
rect 7504 4142 7538 4144
rect 7946 4142 7980 4144
rect 8204 4142 8238 4144
rect 8646 4142 8680 4144
rect 8904 4142 8938 4144
rect 9346 4142 9380 4144
rect 9604 4142 9638 4144
rect 10046 4142 10080 4144
rect 10304 4142 10338 4144
rect -1196 4136 -1162 4138
rect -754 4136 -720 4138
rect -496 4136 -462 4138
rect -54 4136 -20 4138
rect 204 4136 238 4138
rect 646 4136 680 4138
rect 904 4136 938 4138
rect 1346 4136 1380 4138
rect 1604 4136 1638 4138
rect 2046 4136 2080 4138
rect 2304 4136 2338 4138
rect 3746 4136 3780 4138
rect 4004 4136 4038 4138
rect 4446 4136 4480 4138
rect 4704 4136 4738 4138
rect 5146 4136 5180 4138
rect 5404 4136 5438 4138
rect 5846 4136 5880 4138
rect 6104 4136 6138 4138
rect 6546 4136 6580 4138
rect 6804 4136 6838 4138
rect 7246 4136 7280 4138
rect 7504 4136 7538 4138
rect 7946 4136 7980 4138
rect 8204 4136 8238 4138
rect 8646 4136 8680 4138
rect 8904 4136 8938 4138
rect 9346 4136 9380 4138
rect 9604 4136 9638 4138
rect 10046 4136 10080 4138
rect 10304 4136 10338 4138
rect -1196 4108 -1162 4110
rect -754 4108 -720 4110
rect -496 4108 -462 4110
rect -54 4108 -20 4110
rect 204 4108 238 4110
rect 646 4108 680 4110
rect 904 4108 938 4110
rect 1346 4108 1380 4110
rect 1604 4108 1638 4110
rect 2046 4108 2080 4110
rect 2304 4108 2338 4110
rect 3746 4108 3780 4110
rect 4004 4108 4038 4110
rect 4446 4108 4480 4110
rect 4704 4108 4738 4110
rect 5146 4108 5180 4110
rect 5404 4108 5438 4110
rect 5846 4108 5880 4110
rect 6104 4108 6138 4110
rect 6546 4108 6580 4110
rect 6804 4108 6838 4110
rect 7246 4108 7280 4110
rect 7504 4108 7538 4110
rect 7946 4108 7980 4110
rect 8204 4108 8238 4110
rect 8646 4108 8680 4110
rect 8904 4108 8938 4110
rect 9346 4108 9380 4110
rect 9604 4108 9638 4110
rect 10046 4108 10080 4110
rect 10304 4108 10338 4110
rect -1196 4068 -1162 4072
rect -754 4068 -720 4072
rect -496 4068 -462 4072
rect -54 4068 -20 4072
rect 204 4068 238 4072
rect 646 4068 680 4072
rect 904 4068 938 4072
rect 1346 4068 1380 4072
rect 1604 4068 1638 4072
rect 2046 4068 2080 4072
rect 2304 4068 2338 4072
rect 3746 4068 3780 4072
rect 4004 4068 4038 4072
rect 4446 4068 4480 4072
rect 4704 4068 4738 4072
rect 5146 4068 5180 4072
rect 5404 4068 5438 4072
rect 5846 4068 5880 4072
rect 6104 4068 6138 4072
rect 6546 4068 6580 4072
rect 6804 4068 6838 4072
rect 7246 4068 7280 4072
rect 7504 4068 7538 4072
rect 7946 4068 7980 4072
rect 8204 4068 8238 4072
rect 8646 4068 8680 4072
rect 8904 4068 8938 4072
rect 9346 4068 9380 4072
rect 9604 4068 9638 4072
rect 10046 4068 10080 4072
rect 10304 4068 10338 4072
rect -1196 4036 -1162 4038
rect -754 4036 -720 4038
rect -496 4036 -462 4038
rect -54 4036 -20 4038
rect 204 4036 238 4038
rect 646 4036 680 4038
rect 904 4036 938 4038
rect 1346 4036 1380 4038
rect 1604 4036 1638 4038
rect 2046 4036 2080 4038
rect 2304 4036 2338 4038
rect 3746 4036 3780 4038
rect 4004 4036 4038 4038
rect 4446 4036 4480 4038
rect 4704 4036 4738 4038
rect 5146 4036 5180 4038
rect 5404 4036 5438 4038
rect 5846 4036 5880 4038
rect 6104 4036 6138 4038
rect 6546 4036 6580 4038
rect 6804 4036 6838 4038
rect 7246 4036 7280 4038
rect 7504 4036 7538 4038
rect 7946 4036 7980 4038
rect 8204 4036 8238 4038
rect 8646 4036 8680 4038
rect 8904 4036 8938 4038
rect 9346 4036 9380 4038
rect 9604 4036 9638 4038
rect 10046 4036 10080 4038
rect 10304 4036 10338 4038
rect -1196 3998 -1162 4002
rect -754 3998 -720 4002
rect -496 3998 -462 4002
rect -54 3998 -20 4002
rect 204 3998 238 4002
rect 646 3998 680 4002
rect 904 3998 938 4002
rect 1346 3998 1380 4002
rect 1604 3998 1638 4002
rect 2046 3998 2080 4002
rect 2304 3998 2338 4002
rect 3746 3998 3780 4002
rect 4004 3998 4038 4002
rect 4446 3998 4480 4002
rect 4704 3998 4738 4002
rect 5146 3998 5180 4002
rect 5404 3998 5438 4002
rect 5846 3998 5880 4002
rect 6104 3998 6138 4002
rect 6546 3998 6580 4002
rect 6804 3998 6838 4002
rect 7246 3998 7280 4002
rect 7504 3998 7538 4002
rect 7946 3998 7980 4002
rect 8204 3998 8238 4002
rect 8646 3998 8680 4002
rect 8904 3998 8938 4002
rect 9346 3998 9380 4002
rect 9604 3998 9638 4002
rect 10046 3998 10080 4002
rect 10304 3998 10338 4002
rect -1196 3964 -1162 3966
rect -754 3964 -720 3966
rect -496 3964 -462 3966
rect -54 3964 -20 3966
rect 204 3964 238 3966
rect 646 3964 680 3966
rect 904 3964 938 3966
rect 1346 3964 1380 3966
rect 1604 3964 1638 3966
rect 2046 3964 2080 3966
rect 2304 3964 2338 3966
rect 3746 3964 3780 3966
rect 4004 3964 4038 3966
rect 4446 3964 4480 3966
rect 4704 3964 4738 3966
rect 5146 3964 5180 3966
rect 5404 3964 5438 3966
rect 5846 3964 5880 3966
rect 6104 3964 6138 3966
rect 6546 3964 6580 3966
rect 6804 3964 6838 3966
rect 7246 3964 7280 3966
rect 7504 3964 7538 3966
rect 7946 3964 7980 3966
rect 8204 3964 8238 3966
rect 8646 3964 8680 3966
rect 8904 3964 8938 3966
rect 9346 3964 9380 3966
rect 9604 3964 9638 3966
rect 10046 3964 10080 3966
rect 10304 3964 10338 3966
rect -1196 3932 -1162 3934
rect -754 3932 -720 3934
rect -496 3932 -462 3934
rect -54 3932 -20 3934
rect 204 3932 238 3934
rect 646 3932 680 3934
rect 904 3932 938 3934
rect 1346 3932 1380 3934
rect 1604 3932 1638 3934
rect 2046 3932 2080 3934
rect 2304 3932 2338 3934
rect 3746 3932 3780 3934
rect 4004 3932 4038 3934
rect 4446 3932 4480 3934
rect 4704 3932 4738 3934
rect 5146 3932 5180 3934
rect 5404 3932 5438 3934
rect 5846 3932 5880 3934
rect 6104 3932 6138 3934
rect 6546 3932 6580 3934
rect 6804 3932 6838 3934
rect 7246 3932 7280 3934
rect 7504 3932 7538 3934
rect 7946 3932 7980 3934
rect 8204 3932 8238 3934
rect 8646 3932 8680 3934
rect 8904 3932 8938 3934
rect 9346 3932 9380 3934
rect 9604 3932 9638 3934
rect 10046 3932 10080 3934
rect 10304 3932 10338 3934
rect -1196 3926 -1162 3928
rect -754 3926 -720 3928
rect -496 3926 -462 3928
rect -54 3926 -20 3928
rect 204 3926 238 3928
rect 646 3926 680 3928
rect 904 3926 938 3928
rect 1346 3926 1380 3928
rect 1604 3926 1638 3928
rect 2046 3926 2080 3928
rect 2304 3926 2338 3928
rect 3746 3926 3780 3928
rect 4004 3926 4038 3928
rect 4446 3926 4480 3928
rect 4704 3926 4738 3928
rect 5146 3926 5180 3928
rect 5404 3926 5438 3928
rect 5846 3926 5880 3928
rect 6104 3926 6138 3928
rect 6546 3926 6580 3928
rect 6804 3926 6838 3928
rect 7246 3926 7280 3928
rect 7504 3926 7538 3928
rect 7946 3926 7980 3928
rect 8204 3926 8238 3928
rect 8646 3926 8680 3928
rect 8904 3926 8938 3928
rect 9346 3926 9380 3928
rect 9604 3926 9638 3928
rect 10046 3926 10080 3928
rect 10304 3926 10338 3928
rect -1196 3892 -1162 3894
rect -754 3892 -720 3894
rect -496 3892 -462 3894
rect -54 3892 -20 3894
rect 204 3892 238 3894
rect 646 3892 680 3894
rect 904 3892 938 3894
rect 1346 3892 1380 3894
rect 1604 3892 1638 3894
rect 2046 3892 2080 3894
rect 2304 3892 2338 3894
rect 3746 3892 3780 3894
rect 4004 3892 4038 3894
rect 4446 3892 4480 3894
rect 4704 3892 4738 3894
rect 5146 3892 5180 3894
rect 5404 3892 5438 3894
rect 5846 3892 5880 3894
rect 6104 3892 6138 3894
rect 6546 3892 6580 3894
rect 6804 3892 6838 3894
rect 7246 3892 7280 3894
rect 7504 3892 7538 3894
rect 7946 3892 7980 3894
rect 8204 3892 8238 3894
rect 8646 3892 8680 3894
rect 8904 3892 8938 3894
rect 9346 3892 9380 3894
rect 9604 3892 9638 3894
rect 10046 3892 10080 3894
rect 10304 3892 10338 3894
rect -1196 3864 -1162 3866
rect -754 3864 -720 3866
rect -496 3864 -462 3866
rect -54 3864 -20 3866
rect 204 3864 238 3866
rect 646 3864 680 3866
rect 904 3864 938 3866
rect 1346 3864 1380 3866
rect 1604 3864 1638 3866
rect 2046 3864 2080 3866
rect 2304 3864 2338 3866
rect 3746 3864 3780 3866
rect 4004 3864 4038 3866
rect 4446 3864 4480 3866
rect 4704 3864 4738 3866
rect 5146 3864 5180 3866
rect 5404 3864 5438 3866
rect 5846 3864 5880 3866
rect 6104 3864 6138 3866
rect 6546 3864 6580 3866
rect 6804 3864 6838 3866
rect 7246 3864 7280 3866
rect 7504 3864 7538 3866
rect 7946 3864 7980 3866
rect 8204 3864 8238 3866
rect 8646 3864 8680 3866
rect 8904 3864 8938 3866
rect 9346 3864 9380 3866
rect 9604 3864 9638 3866
rect 10046 3864 10080 3866
rect 10304 3864 10338 3866
rect -1196 3854 -1162 3856
rect -754 3854 -720 3856
rect -496 3854 -462 3856
rect -54 3854 -20 3856
rect 204 3854 238 3856
rect 646 3854 680 3856
rect 904 3854 938 3856
rect 1346 3854 1380 3856
rect 1604 3854 1638 3856
rect 2046 3854 2080 3856
rect 2304 3854 2338 3856
rect 3746 3854 3780 3856
rect 4004 3854 4038 3856
rect 4446 3854 4480 3856
rect 4704 3854 4738 3856
rect 5146 3854 5180 3856
rect 5404 3854 5438 3856
rect 5846 3854 5880 3856
rect 6104 3854 6138 3856
rect 6546 3854 6580 3856
rect 6804 3854 6838 3856
rect 7246 3854 7280 3856
rect 7504 3854 7538 3856
rect 7946 3854 7980 3856
rect 8204 3854 8238 3856
rect 8646 3854 8680 3856
rect 8904 3854 8938 3856
rect 9346 3854 9380 3856
rect 9604 3854 9638 3856
rect 10046 3854 10080 3856
rect 10304 3854 10338 3856
rect -1196 3820 -1162 3822
rect -754 3820 -720 3822
rect -496 3820 -462 3822
rect -54 3820 -20 3822
rect 204 3820 238 3822
rect 646 3820 680 3822
rect 904 3820 938 3822
rect 1346 3820 1380 3822
rect 1604 3820 1638 3822
rect 2046 3820 2080 3822
rect 2304 3820 2338 3822
rect 3746 3820 3780 3822
rect 4004 3820 4038 3822
rect 4446 3820 4480 3822
rect 4704 3820 4738 3822
rect 5146 3820 5180 3822
rect 5404 3820 5438 3822
rect 5846 3820 5880 3822
rect 6104 3820 6138 3822
rect 6546 3820 6580 3822
rect 6804 3820 6838 3822
rect 7246 3820 7280 3822
rect 7504 3820 7538 3822
rect 7946 3820 7980 3822
rect 8204 3820 8238 3822
rect 8646 3820 8680 3822
rect 8904 3820 8938 3822
rect 9346 3820 9380 3822
rect 9604 3820 9638 3822
rect 10046 3820 10080 3822
rect 10304 3820 10338 3822
rect -1196 3796 -1162 3798
rect -754 3796 -720 3798
rect -496 3796 -462 3798
rect -54 3796 -20 3798
rect 204 3796 238 3798
rect 646 3796 680 3798
rect 904 3796 938 3798
rect 1346 3796 1380 3798
rect 1604 3796 1638 3798
rect 2046 3796 2080 3798
rect 2304 3796 2338 3798
rect 3746 3796 3780 3798
rect 4004 3796 4038 3798
rect 4446 3796 4480 3798
rect 4704 3796 4738 3798
rect 5146 3796 5180 3798
rect 5404 3796 5438 3798
rect 5846 3796 5880 3798
rect 6104 3796 6138 3798
rect 6546 3796 6580 3798
rect 6804 3796 6838 3798
rect 7246 3796 7280 3798
rect 7504 3796 7538 3798
rect 7946 3796 7980 3798
rect 8204 3796 8238 3798
rect 8646 3796 8680 3798
rect 8904 3796 8938 3798
rect 9346 3796 9380 3798
rect 9604 3796 9638 3798
rect 10046 3796 10080 3798
rect 10304 3796 10338 3798
rect -1196 3782 -1162 3784
rect -754 3782 -720 3784
rect -496 3782 -462 3784
rect -54 3782 -20 3784
rect 204 3782 238 3784
rect 646 3782 680 3784
rect 904 3782 938 3784
rect 1346 3782 1380 3784
rect 1604 3782 1638 3784
rect 2046 3782 2080 3784
rect 2304 3782 2338 3784
rect 3746 3782 3780 3784
rect 4004 3782 4038 3784
rect 4446 3782 4480 3784
rect 4704 3782 4738 3784
rect 5146 3782 5180 3784
rect 5404 3782 5438 3784
rect 5846 3782 5880 3784
rect 6104 3782 6138 3784
rect 6546 3782 6580 3784
rect 6804 3782 6838 3784
rect 7246 3782 7280 3784
rect 7504 3782 7538 3784
rect 7946 3782 7980 3784
rect 8204 3782 8238 3784
rect 8646 3782 8680 3784
rect 8904 3782 8938 3784
rect 9346 3782 9380 3784
rect 9604 3782 9638 3784
rect 10046 3782 10080 3784
rect 10304 3782 10338 3784
rect -1196 3748 -1162 3750
rect -754 3748 -720 3750
rect -496 3748 -462 3750
rect -54 3748 -20 3750
rect 204 3748 238 3750
rect 646 3748 680 3750
rect 904 3748 938 3750
rect 1346 3748 1380 3750
rect 1604 3748 1638 3750
rect 2046 3748 2080 3750
rect 2304 3748 2338 3750
rect 3746 3748 3780 3750
rect 4004 3748 4038 3750
rect 4446 3748 4480 3750
rect 4704 3748 4738 3750
rect 5146 3748 5180 3750
rect 5404 3748 5438 3750
rect 5846 3748 5880 3750
rect 6104 3748 6138 3750
rect 6546 3748 6580 3750
rect 6804 3748 6838 3750
rect 7246 3748 7280 3750
rect 7504 3748 7538 3750
rect 7946 3748 7980 3750
rect 8204 3748 8238 3750
rect 8646 3748 8680 3750
rect 8904 3748 8938 3750
rect 9346 3748 9380 3750
rect 9604 3748 9638 3750
rect 10046 3748 10080 3750
rect 10304 3748 10338 3750
rect -1196 3728 -1162 3730
rect -754 3728 -720 3730
rect -496 3728 -462 3730
rect -54 3728 -20 3730
rect 204 3728 238 3730
rect 646 3728 680 3730
rect 904 3728 938 3730
rect 1346 3728 1380 3730
rect 1604 3728 1638 3730
rect 2046 3728 2080 3730
rect 2304 3728 2338 3730
rect 3746 3728 3780 3730
rect 4004 3728 4038 3730
rect 4446 3728 4480 3730
rect 4704 3728 4738 3730
rect 5146 3728 5180 3730
rect 5404 3728 5438 3730
rect 5846 3728 5880 3730
rect 6104 3728 6138 3730
rect 6546 3728 6580 3730
rect 6804 3728 6838 3730
rect 7246 3728 7280 3730
rect 7504 3728 7538 3730
rect 7946 3728 7980 3730
rect 8204 3728 8238 3730
rect 8646 3728 8680 3730
rect 8904 3728 8938 3730
rect 9346 3728 9380 3730
rect 9604 3728 9638 3730
rect 10046 3728 10080 3730
rect 10304 3728 10338 3730
rect -1196 3710 -1162 3712
rect -754 3710 -720 3712
rect -496 3710 -462 3712
rect -54 3710 -20 3712
rect 204 3710 238 3712
rect 646 3710 680 3712
rect 904 3710 938 3712
rect 1346 3710 1380 3712
rect 1604 3710 1638 3712
rect 2046 3710 2080 3712
rect 2304 3710 2338 3712
rect 3746 3710 3780 3712
rect 4004 3710 4038 3712
rect 4446 3710 4480 3712
rect 4704 3710 4738 3712
rect 5146 3710 5180 3712
rect 5404 3710 5438 3712
rect 5846 3710 5880 3712
rect 6104 3710 6138 3712
rect 6546 3710 6580 3712
rect 6804 3710 6838 3712
rect 7246 3710 7280 3712
rect 7504 3710 7538 3712
rect 7946 3710 7980 3712
rect 8204 3710 8238 3712
rect 8646 3710 8680 3712
rect 8904 3710 8938 3712
rect 9346 3710 9380 3712
rect 9604 3710 9638 3712
rect 10046 3710 10080 3712
rect 10304 3710 10338 3712
rect -1328 3558 -1326 3592
rect -1292 3558 -1288 3592
rect -628 3558 -626 3592
rect -592 3558 -588 3592
rect 72 3558 74 3592
rect 108 3558 112 3592
rect 772 3558 774 3592
rect 808 3558 812 3592
rect 1472 3558 1474 3592
rect 1508 3558 1512 3592
rect 2172 3558 2174 3592
rect 2208 3558 2212 3592
rect 3872 3558 3874 3592
rect 3908 3558 3912 3592
rect 4572 3558 4574 3592
rect 4608 3558 4612 3592
rect 5272 3558 5274 3592
rect 5308 3558 5312 3592
rect 5972 3558 5974 3592
rect 6008 3558 6012 3592
rect 6672 3558 6674 3592
rect 6708 3558 6712 3592
rect 7372 3558 7374 3592
rect 7408 3558 7412 3592
rect 8072 3558 8074 3592
rect 8108 3558 8112 3592
rect 8772 3558 8774 3592
rect 8808 3558 8812 3592
rect 9472 3558 9474 3592
rect 9508 3558 9512 3592
rect 10172 3558 10174 3592
rect 10208 3558 10212 3592
rect 1225 2158 1451 2194
rect 1225 2076 1261 2158
rect 1415 2076 1451 2158
rect 1225 2040 1451 2076
rect 2225 2158 2451 2194
rect 2225 2076 2261 2158
rect 2415 2076 2451 2158
rect 2225 2040 2451 2076
rect 3225 2158 3451 2194
rect 3225 2076 3261 2158
rect 3415 2076 3451 2158
rect 3225 2040 3451 2076
rect 4225 2158 4451 2194
rect 4225 2076 4261 2158
rect 4415 2076 4451 2158
rect 4225 2040 4451 2076
rect 5225 2158 5451 2194
rect 5225 2076 5261 2158
rect 5415 2076 5451 2158
rect 5225 2040 5451 2076
rect 6225 2158 6451 2194
rect 6225 2076 6261 2158
rect 6415 2076 6451 2158
rect 6225 2040 6451 2076
rect 7225 2158 7451 2194
rect 7225 2076 7261 2158
rect 7415 2076 7451 2158
rect 7225 2040 7451 2076
rect 8225 2158 8451 2194
rect 8225 2076 8261 2158
rect 8415 2076 8451 2158
rect 8225 2040 8451 2076
rect 9225 2158 9451 2194
rect 9225 2076 9261 2158
rect 9415 2076 9451 2158
rect 9225 2040 9451 2076
rect 10225 2158 10451 2194
rect 10225 2076 10261 2158
rect 10415 2076 10451 2158
rect 10225 2040 10451 2076
rect 1224 1021 1450 1057
rect 1224 939 1260 1021
rect 1414 939 1450 1021
rect 1224 903 1450 939
rect 2224 1021 2450 1057
rect 2224 939 2260 1021
rect 2414 939 2450 1021
rect 2224 903 2450 939
rect 3224 1021 3450 1057
rect 3224 939 3260 1021
rect 3414 939 3450 1021
rect 3224 903 3450 939
rect 4224 1021 4450 1057
rect 4224 939 4260 1021
rect 4414 939 4450 1021
rect 4224 903 4450 939
rect 5224 1021 5450 1057
rect 5224 939 5260 1021
rect 5414 939 5450 1021
rect 5224 903 5450 939
rect 6224 1021 6450 1057
rect 6224 939 6260 1021
rect 6414 939 6450 1021
rect 6224 903 6450 939
rect 7224 1021 7450 1057
rect 7224 939 7260 1021
rect 7414 939 7450 1021
rect 7224 903 7450 939
rect 8224 1021 8450 1057
rect 8224 939 8260 1021
rect 8414 939 8450 1021
rect 8224 903 8450 939
rect 9224 1021 9450 1057
rect 9224 939 9260 1021
rect 9414 939 9450 1021
rect 9224 903 9450 939
rect 10224 1021 10450 1057
rect 10224 939 10260 1021
rect 10414 939 10450 1021
rect 10224 903 10450 939
<< metal1 >>
rect 1551 8950 1669 9069
rect 2972 8951 4266 9070
rect 4125 7474 4266 8951
rect 4125 7291 11226 7474
rect 2476 6413 2609 6910
rect 2012 6182 2614 6413
rect 3476 6409 3609 6910
rect 3477 6188 3609 6409
rect 12291 3975 12461 5064
rect 12291 3621 13067 3975
rect 2480 2920 4044 3080
rect 956 2287 1083 2411
rect 2586 2397 2711 2920
rect 12291 2520 12461 3621
rect 10711 2397 12461 2520
rect 652 495 852 713
<< metal2 >>
rect 9880 6229 11838 6329
rect -86 5849 60 5951
rect 3845 5849 3991 5951
rect 1786 3404 1937 3492
rect 9752 3405 9920 3493
use contact$4  contact$4_0
timestamp 1635946216
transform 1 0 9996 0 1 6278
box -64 -32 64 32
use diff_pair  diff_pair_0
timestamp 1635946216
transform 1 0 -1557 0 1 3719
box -2909 -799 12037 2621
use current_mirror  current_mirror_0
timestamp 1635946216
transform 1 0 2847 0 1 7379
box -1298 -469 762 1691
use amp  amp_0
timestamp 1635946216
transform 1 0 14597 0 1 6161
box -3371 -1097 4030 1313
use bias_current_mirror  bias_current_mirror_0
timestamp 1635946216
transform 1 0 2122 0 1 3452
box -1470 -2957 8696 488
<< labels >>
flabel metal1 s 1551 8950 1669 9069 2 FreeSans 2000 0 0 0 vdd
port 1 nsew
flabel metal1 s 12747 3625 13063 3972 2 FreeSans 2000 0 0 0 out
port 2 nsew
flabel metal1 s 652 495 852 713 2 FreeSans 2000 0 0 0 vss
port 3 nsew
flabel metal1 s 956 2287 1083 2411 2 FreeSans 2000 0 0 0 bias
port 4 nsew
flabel metal2 s 1786 3404 1937 3492 2 FreeSans 2000 0 0 0 in_n
port 5 nsew
flabel metal2 s 9752 3405 9920 3493 2 FreeSans 2000 0 0 0 in_p
port 6 nsew
flabel metal2 s 3845 5849 3991 5951 2 FreeSans 2000 0 0 0 vss
port 3 nsew
flabel metal2 s -86 5849 60 5951 2 FreeSans 2000 0 0 0 vss
port 3 nsew
<< end >>
