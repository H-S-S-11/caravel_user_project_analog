magic
tech sky130A
magscale 1 2
timestamp 1635946216
<< error_p >>
rect -324 -266 -294 266
rect -258 -200 -228 200
rect 228 -200 258 200
rect 294 -266 324 266
<< nwell >>
rect -294 -576 294 534
<< mvpmos >>
rect -200 -200 200 200
<< mvpdiff >>
rect -258 187 -200 200
rect -258 153 -246 187
rect -212 153 -200 187
rect -258 119 -200 153
rect -258 85 -246 119
rect -212 85 -200 119
rect -258 51 -200 85
rect -258 17 -246 51
rect -212 17 -200 51
rect -258 -17 -200 17
rect -258 -51 -246 -17
rect -212 -51 -200 -17
rect -258 -85 -200 -51
rect -258 -119 -246 -85
rect -212 -119 -200 -85
rect -258 -153 -200 -119
rect -258 -187 -246 -153
rect -212 -187 -200 -153
rect -258 -200 -200 -187
rect 200 187 258 200
rect 200 153 212 187
rect 246 153 258 187
rect 200 119 258 153
rect 200 85 212 119
rect 246 85 258 119
rect 200 51 258 85
rect 200 17 212 51
rect 246 17 258 51
rect 200 -17 258 17
rect 200 -51 212 -17
rect 246 -51 258 -17
rect 200 -85 258 -51
rect 200 -119 212 -85
rect 246 -119 258 -85
rect 200 -153 258 -119
rect 200 -187 212 -153
rect 246 -187 258 -153
rect 200 -200 258 -187
<< mvpdiffc >>
rect -246 153 -212 187
rect -246 85 -212 119
rect -246 17 -212 51
rect -246 -51 -212 -17
rect -246 -119 -212 -85
rect -246 -187 -212 -153
rect 212 153 246 187
rect 212 85 246 119
rect 212 17 246 51
rect 212 -51 246 -17
rect 212 -119 246 -85
rect 212 -187 246 -153
<< poly >>
rect -200 281 200 297
rect -200 247 -153 281
rect -119 247 -85 281
rect -51 247 -17 281
rect 17 247 51 281
rect 85 247 119 281
rect 153 247 200 281
rect -200 200 200 247
rect -200 -247 200 -200
rect -200 -281 -153 -247
rect -119 -281 -85 -247
rect -51 -281 -17 -247
rect 17 -281 51 -247
rect 85 -281 119 -247
rect 153 -281 200 -247
rect -200 -297 200 -281
<< polycont >>
rect -153 247 -119 281
rect -85 247 -51 281
rect -17 247 17 281
rect 51 247 85 281
rect 119 247 153 281
rect -153 -281 -119 -247
rect -85 -281 -51 -247
rect -17 -281 17 -247
rect 51 -281 85 -247
rect 119 -281 153 -247
<< locali >>
rect -200 247 -161 281
rect -119 247 -89 281
rect -51 247 -17 281
rect 17 247 51 281
rect 89 247 119 281
rect 161 247 200 281
rect -246 187 -212 204
rect -246 119 -212 127
rect -246 51 -212 55
rect -246 -55 -212 -51
rect -246 -127 -212 -119
rect -246 -204 -212 -187
rect 212 187 246 204
rect 212 119 246 127
rect 212 51 246 55
rect 212 -55 246 -51
rect 212 -127 246 -119
rect 212 -204 246 -187
rect -200 -281 -161 -247
rect -119 -281 -89 -247
rect -51 -281 -17 -247
rect 17 -281 51 -247
rect 89 -281 119 -247
rect 161 -281 200 -247
<< viali >>
rect -161 247 -153 281
rect -153 247 -127 281
rect -89 247 -85 281
rect -85 247 -55 281
rect -17 247 17 281
rect 55 247 85 281
rect 85 247 89 281
rect 127 247 153 281
rect 153 247 161 281
rect -246 153 -212 161
rect -246 127 -212 153
rect -246 85 -212 89
rect -246 55 -212 85
rect -246 -17 -212 17
rect -246 -85 -212 -55
rect -246 -89 -212 -85
rect -246 -153 -212 -127
rect -246 -161 -212 -153
rect 212 153 246 161
rect 212 127 246 153
rect 212 85 246 89
rect 212 55 246 85
rect 212 -17 246 17
rect 212 -85 246 -55
rect 212 -89 246 -85
rect 212 -153 246 -127
rect 212 -161 246 -153
rect -161 -281 -153 -247
rect -153 -281 -127 -247
rect -89 -281 -85 -247
rect -85 -281 -55 -247
rect -17 -281 17 -247
rect 55 -281 85 -247
rect 85 -281 89 -247
rect 127 -281 153 -247
rect 153 -281 161 -247
<< metal1 >>
rect -196 281 196 287
rect -196 247 -161 281
rect -127 247 -89 281
rect -55 247 -17 281
rect 17 247 55 281
rect 89 247 127 281
rect 161 247 196 281
rect -196 241 196 247
rect -252 161 -206 200
rect -252 127 -246 161
rect -212 127 -206 161
rect -252 89 -206 127
rect -252 55 -246 89
rect -212 55 -206 89
rect -252 17 -206 55
rect -252 -17 -246 17
rect -212 -17 -206 17
rect -252 -55 -206 -17
rect -252 -89 -246 -55
rect -212 -89 -206 -55
rect -252 -127 -206 -89
rect -252 -161 -246 -127
rect -212 -161 -206 -127
rect -252 -200 -206 -161
rect 206 161 252 200
rect 206 127 212 161
rect 246 127 252 161
rect 206 89 252 127
rect 206 55 212 89
rect 246 55 252 89
rect 206 17 252 55
rect 206 -17 212 17
rect 246 -17 252 17
rect 206 -55 252 -17
rect 206 -89 212 -55
rect 246 -89 252 -55
rect 206 -127 252 -89
rect 206 -161 212 -127
rect 246 -161 252 -127
rect 206 -200 252 -161
rect -196 -247 196 -241
rect -196 -281 -161 -247
rect -127 -281 -89 -247
rect -55 -281 -17 -247
rect 17 -281 55 -247
rect 89 -281 127 -247
rect 161 -281 196 -247
rect -196 -287 196 -281
<< end >>
