magic
tech sky130A
timestamp 1633983039
<< dnwell >>
rect -791 -371 409 429
<< nwell >>
rect -751 -271 -531 329
<< pwell >>
rect -461 329 -341 429
rect -311 329 -251 429
rect -491 -271 309 329
<< nmos >>
rect -211 59 -193 159
rect 189 59 207 159
rect -211 -151 -193 -51
rect 189 -151 207 -51
<< nsonos >>
rect -82 55 -64 155
rect -33 55 -15 155
rect 16 55 34 155
rect 65 55 83 155
rect -82 -156 -64 -56
rect -33 -156 -15 -56
rect 16 -156 34 -56
rect 65 -156 83 -56
<< ndiff >>
rect -251 149 -211 159
rect -251 69 -241 149
rect -221 69 -211 149
rect -251 59 -211 69
rect -193 149 -151 159
rect -193 69 -181 149
rect -161 69 -151 149
rect -193 59 -151 69
rect -112 149 -82 155
rect -112 61 -106 149
rect -88 61 -82 149
rect -112 55 -82 61
rect -64 55 -33 155
rect -15 55 16 155
rect 34 55 65 155
rect 83 149 113 155
rect 83 61 89 149
rect 107 61 113 149
rect 83 55 113 61
rect 149 149 189 159
rect 149 69 159 149
rect 179 69 189 149
rect 149 59 189 69
rect 207 149 249 159
rect 207 69 219 149
rect 239 69 249 149
rect 207 59 249 69
rect -251 -61 -211 -51
rect -251 -141 -241 -61
rect -221 -141 -211 -61
rect -251 -151 -211 -141
rect -193 -61 -151 -51
rect -193 -141 -181 -61
rect -161 -141 -151 -61
rect -193 -151 -151 -141
rect -112 -62 -82 -56
rect -112 -150 -106 -62
rect -88 -150 -82 -62
rect -112 -156 -82 -150
rect -64 -156 -33 -56
rect -15 -156 16 -56
rect 34 -156 65 -56
rect 83 -62 113 -56
rect 83 -150 89 -62
rect 107 -150 113 -62
rect 83 -156 113 -150
rect 149 -61 189 -51
rect 149 -141 159 -61
rect 179 -141 189 -61
rect 149 -151 189 -141
rect 207 -61 249 -51
rect 207 -141 219 -61
rect 239 -141 249 -61
rect 207 -151 249 -141
<< ndiffc >>
rect -241 69 -221 149
rect -181 69 -161 149
rect -106 61 -88 149
rect 89 61 107 149
rect 159 69 179 149
rect 219 69 239 149
rect -241 -141 -221 -61
rect -181 -141 -161 -61
rect -106 -150 -88 -62
rect 89 -150 107 -62
rect 159 -141 179 -61
rect 219 -141 239 -61
<< psubdiff >>
rect -461 139 -341 159
rect -461 -131 -441 139
rect -361 -131 -341 139
rect -461 -151 -341 -131
<< nsubdiff >>
rect -731 289 -551 309
rect -731 -231 -711 289
rect -571 -231 -551 289
rect -731 -251 -551 -231
<< psubdiffcont >>
rect -441 -131 -361 139
<< nsubdiffcont >>
rect -711 -231 -571 289
<< poly >>
rect -36 279 -6 289
rect -36 259 -31 279
rect -11 259 -6 279
rect -36 249 -6 259
rect 64 279 94 289
rect 64 259 69 279
rect 89 259 94 279
rect 64 249 94 259
rect -221 219 -181 229
rect -221 199 -211 219
rect -191 199 -181 219
rect -221 189 -181 199
rect -96 219 -61 229
rect -96 199 -91 219
rect -71 199 -61 219
rect -96 189 -61 199
rect -211 159 -193 189
rect -82 155 -64 189
rect -33 155 -15 249
rect 14 219 44 229
rect 14 199 19 219
rect 39 199 44 219
rect 14 189 44 199
rect 16 155 34 189
rect 65 155 83 249
rect 179 219 219 229
rect 179 199 189 219
rect 209 199 219 219
rect 179 189 219 199
rect 189 159 207 189
rect -211 -51 -193 59
rect -82 -56 -64 55
rect -33 -56 -15 55
rect 16 -56 34 55
rect 65 -56 83 55
rect 189 -51 207 59
rect -211 -171 -193 -151
rect -82 -171 -64 -156
rect -33 -171 -15 -156
rect 16 -171 34 -156
rect 65 -171 83 -156
rect 189 -171 207 -151
<< polycont >>
rect -31 259 -11 279
rect 69 259 89 279
rect -211 199 -191 219
rect -91 199 -71 219
rect 19 199 39 219
rect 189 199 209 219
<< locali >>
rect -731 289 -551 429
rect -731 -231 -711 289
rect -571 -231 -551 289
rect -461 139 -341 429
rect -461 -131 -441 139
rect -361 -131 -341 139
rect -461 -151 -341 -131
rect -311 159 -251 429
rect -221 219 -181 429
rect -141 359 -111 429
rect -141 329 -61 359
rect -221 199 -211 219
rect -191 199 -181 219
rect -221 189 -181 199
rect -96 219 -61 329
rect -36 279 -6 429
rect -36 259 -31 279
rect -11 259 -6 279
rect -36 249 -6 259
rect -96 199 -91 219
rect -71 199 -61 219
rect -96 189 -61 199
rect 14 219 44 429
rect 109 359 139 429
rect 64 329 139 359
rect 64 279 94 329
rect 64 259 69 279
rect 89 259 94 279
rect 64 249 94 259
rect 14 199 19 219
rect 39 199 44 219
rect 14 189 44 199
rect 179 219 219 429
rect 179 199 189 219
rect 209 199 219 219
rect 179 189 219 199
rect -311 149 -221 159
rect -311 69 -241 149
rect -311 59 -221 69
rect -181 149 -151 159
rect -106 149 -88 157
rect -161 69 -106 149
rect -181 61 -106 69
rect -181 59 -88 61
rect -311 -51 -251 59
rect -106 53 -88 59
rect 89 149 107 157
rect 149 149 179 159
rect 107 69 159 149
rect 107 61 179 69
rect 89 59 179 61
rect 219 149 409 159
rect 239 69 409 149
rect 219 59 409 69
rect 89 53 107 59
rect -311 -61 -221 -51
rect -311 -141 -241 -61
rect -311 -151 -221 -141
rect -181 -61 -151 -51
rect -106 -61 -88 -54
rect -161 -62 -88 -61
rect -161 -141 -106 -62
rect -181 -150 -106 -141
rect -181 -151 -88 -150
rect -106 -158 -88 -151
rect 89 -61 107 -54
rect 149 -61 179 -51
rect 89 -62 159 -61
rect 107 -141 159 -62
rect 107 -150 179 -141
rect 89 -151 179 -150
rect 219 -61 409 -51
rect 239 -141 409 -61
rect 219 -151 409 -141
rect 89 -158 107 -151
rect -731 -251 -551 -231
<< properties >>
string gencell sky130_fd_bs_flash__special_sonosfet_star
string parameters w 1 l 0.18 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
