magic
tech sky130A
timestamp 1634764606
<< nwell >>
rect 800 -600 2150 900
<< pwell >>
rect -400 -600 650 900
<< nnmos >>
rect 400 -500 450 500
<< mvpmos >>
rect 1000 -500 1050 200
rect 1200 -500 1250 200
<< mvndiff >>
rect 300 490 400 500
rect 300 -490 310 490
rect 380 -490 400 490
rect 300 -500 400 -490
rect 450 490 550 500
rect 450 -490 470 490
rect 540 -490 550 490
rect 450 -500 550 -490
<< mvpdiff >>
rect 900 190 1000 200
rect 900 -490 910 190
rect 980 -490 1000 190
rect 900 -500 1000 -490
rect 1050 180 1200 200
rect 1050 -490 1070 180
rect 1180 -490 1200 180
rect 1050 -500 1200 -490
rect 1250 190 1350 200
rect 1250 -490 1270 190
rect 1340 -490 1350 190
rect 1250 -500 1350 -490
<< mvndiffc >>
rect 310 -490 380 490
rect 470 -490 540 490
<< mvpdiffc >>
rect 910 -490 980 190
rect 1070 -490 1180 180
rect 1270 -490 1340 190
<< mvpsubdiff >>
rect -400 850 100 900
rect -400 450 -350 850
rect 50 450 100 850
rect -400 400 100 450
<< mvnsubdiff >>
rect 1650 -50 2100 0
rect 1650 -450 1700 -50
rect 2050 -450 2100 -50
rect 1650 -500 2100 -450
<< mvpsubdiffcont >>
rect -350 450 50 850
<< mvnsubdiffcont >>
rect 1700 -450 2050 -50
<< poly >>
rect 300 650 550 700
rect 300 600 350 650
rect 500 600 550 650
rect 300 550 550 600
rect 400 500 450 550
rect 1000 350 1250 400
rect 1000 300 1050 350
rect 1200 300 1250 350
rect 1000 250 1250 300
rect 1000 200 1050 250
rect 1200 200 1250 250
rect 400 -550 450 -500
rect 1000 -550 1050 -500
rect 1200 -550 1250 -500
rect 300 -600 550 -550
rect 300 -650 350 -600
rect 500 -650 550 -600
rect 300 -700 550 -650
rect 1000 -600 1250 -550
rect 1000 -650 1050 -600
rect 1200 -650 1250 -600
rect 1000 -700 1250 -650
<< polycont >>
rect 350 600 500 650
rect 1050 300 1200 350
rect 350 -650 500 -600
rect 1050 -650 1200 -600
<< locali >>
rect -400 850 100 900
rect -400 450 -350 850
rect 50 450 100 850
rect 300 650 550 1100
rect 300 600 350 650
rect 500 600 550 650
rect 300 550 550 600
rect -400 400 100 450
rect 470 490 900 500
rect 540 480 900 490
rect 540 170 570 480
rect 880 200 900 480
rect 1000 350 1250 1100
rect 1000 300 1050 350
rect 1200 300 1250 350
rect 1000 250 1250 300
rect 880 190 980 200
rect 880 170 910 190
rect 540 -490 910 170
rect 470 -500 980 -490
rect 1270 190 1350 200
rect 1340 -490 1350 190
rect 1270 -500 1350 -490
rect 1650 -50 2150 0
rect 1650 -450 1700 -50
rect 2100 -450 2150 -50
rect 1650 -500 2150 -450
rect 300 -600 550 -550
rect 300 -650 350 -600
rect 500 -650 550 -600
rect 300 -750 550 -650
rect 1000 -600 1250 -550
rect 1000 -650 1050 -600
rect 1200 -650 1250 -600
rect 1000 -750 1250 -650
<< viali >>
rect -350 450 50 850
rect 220 490 380 500
rect 220 -490 310 490
rect 310 -490 380 490
rect 220 -500 380 -490
rect 570 170 880 480
rect 1070 180 1180 200
rect 1070 -490 1180 180
rect 1070 -500 1180 -490
rect 1350 -500 1500 500
rect 1700 -450 2050 -50
rect 2050 -450 2100 -50
<< metal1 >>
rect -400 850 100 900
rect -400 450 -350 850
rect 50 450 100 850
rect -400 400 100 450
rect 200 500 400 520
rect 200 0 220 500
rect -500 -400 220 0
rect 200 -500 220 -400
rect 380 0 400 500
rect 550 500 2250 800
rect 550 480 1350 500
rect 550 170 570 480
rect 880 300 1350 480
rect 880 170 900 300
rect 550 150 900 170
rect 1050 200 1200 210
rect 1050 0 1070 200
rect 380 -400 1070 0
rect 380 -500 400 -400
rect 200 -520 400 -500
rect 1050 -500 1070 -400
rect 1180 -500 1200 200
rect 1050 -520 1200 -500
rect 1330 -500 1350 300
rect 1500 400 2250 500
rect 1500 -500 1520 400
rect 1650 -50 2150 0
rect 1650 -450 1700 -50
rect 2100 -450 2150 -50
rect 1650 -500 2150 -450
rect 1330 -520 1520 -500
<< via1 >>
rect -350 450 50 850
rect 1700 -450 2100 -50
<< metal2 >>
rect -400 850 100 1100
rect -400 450 -350 850
rect 50 450 100 850
rect -400 -750 100 450
rect 1650 -50 2150 1100
rect 1650 -450 1700 -50
rect 2100 -450 2150 -50
rect 1650 -750 2150 -450
<< labels >>
rlabel metal1 2200 400 2250 800 1 VOUT
port 1 n
rlabel metal1 -500 -400 -450 0 1 VIN
port 2 n
rlabel locali 300 1050 550 1100 1 EN
port 3 n
rlabel locali 1000 1050 1250 1100 1 ENB
port 4 n
rlabel metal2 1650 1050 2150 1100 1 VDD3v3
port 5 n
rlabel metal2 -400 1050 100 1100 1 VGND
port 6 n
rlabel metal2 -400 -750 100 -700 1 VGND
port 6 n
rlabel metal2 1650 -750 2150 -700 1 VDD3v3
port 5 n
rlabel locali 300 -750 550 -700 1 EN
port 3 n
rlabel locali 1000 -750 1250 -700 1 ENB
port 4 n
<< end >>
