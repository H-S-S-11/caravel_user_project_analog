magic
tech sky130A
timestamp 1635946216
<< end >>
