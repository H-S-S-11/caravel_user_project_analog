magic
tech sky130A
magscale 1 2
timestamp 1632244313
<< pwell >>
rect -377 -776 377 776
<< nnmos >>
rect -149 318 -29 518
rect 29 318 149 518
rect -149 -100 -29 100
rect 29 -100 149 100
rect -149 -518 -29 -318
rect 29 -518 149 -318
<< mvndiff >>
rect -207 506 -149 518
rect -207 330 -195 506
rect -161 330 -149 506
rect -207 318 -149 330
rect -29 506 29 518
rect -29 330 -17 506
rect 17 330 29 506
rect -29 318 29 330
rect 149 506 207 518
rect 149 330 161 506
rect 195 330 207 506
rect 149 318 207 330
rect -207 88 -149 100
rect -207 -88 -195 88
rect -161 -88 -149 88
rect -207 -100 -149 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 149 88 207 100
rect 149 -88 161 88
rect 195 -88 207 88
rect 149 -100 207 -88
rect -207 -330 -149 -318
rect -207 -506 -195 -330
rect -161 -506 -149 -330
rect -207 -518 -149 -506
rect -29 -330 29 -318
rect -29 -506 -17 -330
rect 17 -506 29 -330
rect -29 -518 29 -506
rect 149 -330 207 -318
rect 149 -506 161 -330
rect 195 -506 207 -330
rect 149 -518 207 -506
<< mvndiffc >>
rect -195 330 -161 506
rect -17 330 17 506
rect 161 330 195 506
rect -195 -88 -161 88
rect -17 -88 17 88
rect 161 -88 195 88
rect -195 -506 -161 -330
rect -17 -506 17 -330
rect 161 -506 195 -330
<< mvpsubdiff >>
rect -341 728 341 740
rect -341 694 -233 728
rect 233 694 341 728
rect -341 682 341 694
rect -341 632 -283 682
rect -341 -632 -329 632
rect -295 -632 -283 632
rect 283 632 341 682
rect -341 -682 -283 -632
rect 283 -632 295 632
rect 329 -632 341 632
rect 283 -682 341 -632
rect -341 -694 341 -682
rect -341 -728 -233 -694
rect 233 -728 341 -694
rect -341 -740 341 -728
<< mvpsubdiffcont >>
rect -233 694 233 728
rect -329 -632 -295 632
rect 295 -632 329 632
rect -233 -728 233 -694
<< poly >>
rect -149 590 -29 606
rect -149 556 -133 590
rect -45 556 -29 590
rect -149 518 -29 556
rect 29 590 149 606
rect 29 556 45 590
rect 133 556 149 590
rect 29 518 149 556
rect -149 280 -29 318
rect -149 246 -133 280
rect -45 246 -29 280
rect -149 230 -29 246
rect 29 280 149 318
rect 29 246 45 280
rect 133 246 149 280
rect 29 230 149 246
rect -149 172 -29 188
rect -149 138 -133 172
rect -45 138 -29 172
rect -149 100 -29 138
rect 29 172 149 188
rect 29 138 45 172
rect 133 138 149 172
rect 29 100 149 138
rect -149 -138 -29 -100
rect -149 -172 -133 -138
rect -45 -172 -29 -138
rect -149 -188 -29 -172
rect 29 -138 149 -100
rect 29 -172 45 -138
rect 133 -172 149 -138
rect 29 -188 149 -172
rect -149 -246 -29 -230
rect -149 -280 -133 -246
rect -45 -280 -29 -246
rect -149 -318 -29 -280
rect 29 -246 149 -230
rect 29 -280 45 -246
rect 133 -280 149 -246
rect 29 -318 149 -280
rect -149 -556 -29 -518
rect -149 -590 -133 -556
rect -45 -590 -29 -556
rect -149 -606 -29 -590
rect 29 -556 149 -518
rect 29 -590 45 -556
rect 133 -590 149 -556
rect 29 -606 149 -590
<< polycont >>
rect -133 556 -45 590
rect 45 556 133 590
rect -133 246 -45 280
rect 45 246 133 280
rect -133 138 -45 172
rect 45 138 133 172
rect -133 -172 -45 -138
rect 45 -172 133 -138
rect -133 -280 -45 -246
rect 45 -280 133 -246
rect -133 -590 -45 -556
rect 45 -590 133 -556
<< locali >>
rect -329 694 -233 728
rect 233 694 329 728
rect -329 632 -295 694
rect 295 632 329 694
rect -149 556 -133 590
rect -45 556 -29 590
rect 29 556 45 590
rect 133 556 149 590
rect -195 506 -161 522
rect -195 314 -161 330
rect -17 506 17 522
rect -17 314 17 330
rect 161 506 195 522
rect 161 314 195 330
rect -149 246 -133 280
rect -45 246 -29 280
rect 29 246 45 280
rect 133 246 149 280
rect -149 138 -133 172
rect -45 138 -29 172
rect 29 138 45 172
rect 133 138 149 172
rect -195 88 -161 104
rect -195 -104 -161 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 161 88 195 104
rect 161 -104 195 -88
rect -149 -172 -133 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 133 -172 149 -138
rect -149 -280 -133 -246
rect -45 -280 -29 -246
rect 29 -280 45 -246
rect 133 -280 149 -246
rect -195 -330 -161 -314
rect -195 -522 -161 -506
rect -17 -330 17 -314
rect -17 -522 17 -506
rect 161 -330 195 -314
rect 161 -522 195 -506
rect -149 -590 -133 -556
rect -45 -590 -29 -556
rect 29 -590 45 -556
rect 133 -590 149 -556
rect -329 -694 -295 -632
rect 295 -694 329 -632
rect -329 -728 -233 -694
rect 233 -728 329 -694
<< properties >>
string gencell sky130_fd_pr__nfet_03v3_nvt
string FIXED_BBOX -312 -711 312 711
string parameters w 1 l 0.6 m 3 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
