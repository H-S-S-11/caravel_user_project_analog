magic
tech sky130A
magscale 1 2
timestamp 1632393576
<< nwell >>
rect -214 -1773 214 1773
<< pmos >>
rect -18 954 18 1554
rect -18 118 18 718
rect -18 -718 18 -118
rect -18 -1554 18 -954
<< pdiff >>
rect -76 1542 -18 1554
rect -76 966 -64 1542
rect -30 966 -18 1542
rect -76 954 -18 966
rect 18 1542 76 1554
rect 18 966 30 1542
rect 64 966 76 1542
rect 18 954 76 966
rect -76 706 -18 718
rect -76 130 -64 706
rect -30 130 -18 706
rect -76 118 -18 130
rect 18 706 76 718
rect 18 130 30 706
rect 64 130 76 706
rect 18 118 76 130
rect -76 -130 -18 -118
rect -76 -706 -64 -130
rect -30 -706 -18 -130
rect -76 -718 -18 -706
rect 18 -130 76 -118
rect 18 -706 30 -130
rect 64 -706 76 -130
rect 18 -718 76 -706
rect -76 -966 -18 -954
rect -76 -1542 -64 -966
rect -30 -1542 -18 -966
rect -76 -1554 -18 -1542
rect 18 -966 76 -954
rect 18 -1542 30 -966
rect 64 -1542 76 -966
rect 18 -1554 76 -1542
<< pdiffc >>
rect -64 966 -30 1542
rect 30 966 64 1542
rect -64 130 -30 706
rect 30 130 64 706
rect -64 -706 -30 -130
rect 30 -706 64 -130
rect -64 -1542 -30 -966
rect 30 -1542 64 -966
<< nsubdiff >>
rect -178 1703 -82 1737
rect 82 1703 178 1737
rect -178 1641 -144 1703
rect 144 1641 178 1703
rect -178 -1703 -144 -1641
rect 144 -1703 178 -1641
rect -178 -1737 -82 -1703
rect 82 -1737 178 -1703
<< nsubdiffcont >>
rect -82 1703 82 1737
rect -178 -1641 -144 1641
rect 144 -1641 178 1641
rect -82 -1737 82 -1703
<< poly >>
rect -33 1635 33 1651
rect -33 1601 -17 1635
rect 17 1601 33 1635
rect -33 1585 33 1601
rect -18 1554 18 1585
rect -18 923 18 954
rect -33 907 33 923
rect -33 873 -17 907
rect 17 873 33 907
rect -33 857 33 873
rect -33 799 33 815
rect -33 765 -17 799
rect 17 765 33 799
rect -33 749 33 765
rect -18 718 18 749
rect -18 87 18 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -18 -118 18 -87
rect -18 -749 18 -718
rect -33 -765 33 -749
rect -33 -799 -17 -765
rect 17 -799 33 -765
rect -33 -815 33 -799
rect -33 -873 33 -857
rect -33 -907 -17 -873
rect 17 -907 33 -873
rect -33 -923 33 -907
rect -18 -954 18 -923
rect -18 -1585 18 -1554
rect -33 -1601 33 -1585
rect -33 -1635 -17 -1601
rect 17 -1635 33 -1601
rect -33 -1651 33 -1635
<< polycont >>
rect -17 1601 17 1635
rect -17 873 17 907
rect -17 765 17 799
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -799 17 -765
rect -17 -907 17 -873
rect -17 -1635 17 -1601
<< locali >>
rect -178 1703 -82 1737
rect 82 1703 178 1737
rect -178 1641 -144 1703
rect 144 1641 178 1703
rect -33 1601 -17 1635
rect 17 1601 33 1635
rect -64 1542 -30 1558
rect -64 950 -30 966
rect 30 1542 64 1558
rect 30 950 64 966
rect -33 873 -17 907
rect 17 873 33 907
rect -33 765 -17 799
rect 17 765 33 799
rect -64 706 -30 722
rect -64 114 -30 130
rect 30 706 64 722
rect 30 114 64 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -64 -130 -30 -114
rect -64 -722 -30 -706
rect 30 -130 64 -114
rect 30 -722 64 -706
rect -33 -799 -17 -765
rect 17 -799 33 -765
rect -33 -907 -17 -873
rect 17 -907 33 -873
rect -64 -966 -30 -950
rect -64 -1558 -30 -1542
rect 30 -966 64 -950
rect 30 -1558 64 -1542
rect -33 -1635 -17 -1601
rect 17 -1635 33 -1601
rect -178 -1703 -144 -1641
rect 144 -1703 178 -1641
rect -178 -1737 -82 -1703
rect 82 -1737 178 -1703
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -161 -1720 161 1720
string parameters w 3 l 0.18 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
