* scale: 1e6 units = 1 micron

* This is a 1.8V version: make sure expected inputs in range

.subckt comparator-diffamp VOP VON VOUT VGND VPWR

*load transistors
X0 VPWR VONAMP VOPAMP VPWR sky130_fd_pr__pfet_01v8 w=3e+06u l=0.18e+6u
X1 VPWR VONAMP VONAMP VPWR sky130_fd_pr__pfet_01v8 w=3e+06u l=0.18e+6u

*diff pair
X2 VOPAMP VOP ISINK VGND sky130_fd_pr__nfet_01v8 w=1e+06u l=0.18e+6u
X3 VONAMP VON ISINK VGND sky130_fd_pr__nfet_01v8 w=1e+06u l=0.18e+6u

* current source
X4 ISINK VONAMP VGND VGND sky130_fd_pr__nfet_01v8 w=1e+06u l=0.18e+6u

*output inverter
X5 VPWR VOPAMP VOUT VPWR sky130_fd_pr__pfet_01v8 w=2e+06u l=0.15e+6u
X6 VOUT VOPAMP VGND VGND sky130_fd_pr__nfet_01v8 w=1e+06u l=0.15e+6u


.ends