magic
tech sky130A
timestamp 1636296152
<< locali >>
rect 1076 4352 1145 4385
rect 1576 4352 1645 4385
rect 989 4053 1006 4257
rect 1489 4053 1506 4257
rect 989 3683 1006 3887
rect 1489 3683 1506 3887
rect 10541 3740 10574 3810
rect 1074 3550 1143 3583
rect 1574 3550 1643 3583
rect 5935 3522 6004 3555
rect 6385 3522 6454 3555
rect 6835 3522 6904 3555
rect 7285 3522 7354 3555
rect 7735 3522 7804 3555
rect 8185 3522 8254 3555
rect 8635 3522 8704 3555
rect 9085 3522 9154 3555
rect 5848 3223 5865 3427
rect 6077 3223 6094 3427
rect 6298 3223 6315 3427
rect 6527 3223 6544 3427
rect 6748 3223 6765 3427
rect 6977 3223 6994 3427
rect 7198 3223 7215 3427
rect 7427 3223 7444 3427
rect 7648 3223 7665 3427
rect 7877 3223 7894 3427
rect 8098 3223 8115 3427
rect 8327 3223 8344 3427
rect 8548 3223 8565 3427
rect 8777 3223 8794 3427
rect 8998 3223 9015 3427
rect 9227 3223 9244 3427
rect 5848 2853 5865 3057
rect 6077 2853 6094 3057
rect 6298 2853 6315 3057
rect 6527 2853 6544 3057
rect 6748 2853 6765 3057
rect 6977 2853 6994 3057
rect 7198 2853 7215 3057
rect 7427 2853 7444 3057
rect 7648 2853 7665 3057
rect 7877 2853 7894 3057
rect 8098 2853 8115 3057
rect 8327 2853 8344 3057
rect 8548 2853 8565 3057
rect 8777 2853 8794 3057
rect 8998 2853 9015 3057
rect 9227 2853 9244 3057
rect 10720 3028 10789 3244
rect -2104 2834 -2004 2851
rect -1754 2834 -1654 2851
rect -1404 2834 -1304 2851
rect -1054 2834 -954 2851
rect -704 2834 -604 2851
rect -354 2834 -254 2851
rect -4 2834 96 2851
rect 346 2834 446 2851
rect 696 2834 796 2851
rect 1046 2834 1146 2851
rect 1896 2834 1996 2851
rect 2246 2834 2346 2851
rect 2596 2834 2696 2851
rect 2946 2834 3046 2851
rect 3296 2834 3396 2851
rect 3646 2834 3746 2851
rect 3996 2834 4096 2851
rect 4346 2834 4446 2851
rect 4696 2834 4796 2851
rect 5046 2834 5146 2851
rect 5933 2720 6002 2753
rect 6383 2720 6452 2753
rect 6833 2720 6902 2753
rect 7283 2720 7352 2753
rect 7733 2720 7802 2753
rect 8183 2720 8252 2753
rect 8633 2720 8702 2753
rect 9083 2720 9152 2753
rect -2104 1779 -2004 1796
rect -1754 1779 -1654 1796
rect -1404 1779 -1304 1796
rect -1054 1779 -954 1796
rect -704 1779 -604 1796
rect -354 1779 -254 1796
rect -4 1779 96 1796
rect 346 1779 446 1796
rect 696 1779 796 1796
rect 1046 1779 1146 1796
rect 1896 1779 1996 1796
rect 2246 1779 2346 1796
rect 2596 1779 2696 1796
rect 2946 1779 3046 1796
rect 3296 1779 3396 1796
rect 3646 1779 3746 1796
rect 3996 1779 4096 1796
rect 4346 1779 4446 1796
rect 4696 1779 4796 1796
rect 5046 1779 5146 1796
rect 635 1042 704 1075
rect 1135 1042 1204 1075
rect 1635 1042 1704 1075
rect 2135 1042 2204 1075
rect 2635 1042 2704 1075
rect 3135 1042 3204 1075
rect 3635 1042 3704 1075
rect 4135 1042 4204 1075
rect 4635 1042 4704 1075
rect 5135 1042 5204 1075
rect 567 977 767 994
rect 1067 977 1267 994
rect 1567 977 1767 994
rect 2067 977 2267 994
rect 2567 977 2767 994
rect 3067 977 3267 994
rect 3567 977 3767 994
rect 4067 977 4267 994
rect 4567 977 4767 994
rect 5067 977 5267 994
rect 544 856 561 960
rect 773 856 790 960
rect 1044 856 1061 960
rect 1544 856 1561 960
rect 1773 856 1790 960
rect 2044 856 2061 960
rect 2273 856 2290 960
rect 2544 856 2561 960
rect 2773 856 2790 960
rect 3044 856 3061 960
rect 3273 856 3290 960
rect 3544 856 3561 960
rect 3773 856 3790 960
rect 4044 856 4061 960
rect 4273 856 4290 960
rect 4544 856 4561 960
rect 4773 856 4790 960
rect 5044 856 5061 960
rect 5273 856 5290 960
rect 567 822 767 839
rect 1067 822 1267 839
rect 1567 822 1767 839
rect 2067 822 2267 839
rect 2567 822 2767 839
rect 3067 822 3267 839
rect 3567 822 3767 839
rect 4067 822 4267 839
rect 4567 822 4767 839
rect 5067 822 5267 839
rect 567 727 767 744
rect 1067 727 1267 744
rect 1567 727 1767 744
rect 2067 727 2267 744
rect 2567 727 2767 744
rect 3067 727 3267 744
rect 3567 727 3767 744
rect 4067 727 4267 744
rect 4567 727 4767 744
rect 5067 727 5267 744
rect 544 606 561 710
rect 773 606 790 710
rect 1044 606 1061 710
rect 1544 606 1561 710
rect 1773 606 1790 710
rect 2044 606 2061 710
rect 2273 606 2290 710
rect 2544 606 2561 710
rect 2773 606 2790 710
rect 3044 606 3061 710
rect 3273 606 3290 710
rect 3544 606 3561 710
rect 3773 606 3790 710
rect 4044 606 4061 710
rect 4273 606 4290 710
rect 4544 606 4561 710
rect 4773 606 4790 710
rect 5044 606 5061 710
rect 5273 606 5290 710
rect 567 572 767 589
rect 1067 572 1267 589
rect 1567 572 1767 589
rect 2067 572 2267 589
rect 2567 572 2767 589
rect 3067 572 3267 589
rect 3567 572 3767 589
rect 4067 572 4267 589
rect 4567 572 4767 589
rect 5067 572 5267 589
rect 634 474 703 507
rect 1134 474 1203 507
rect 1634 474 1703 507
rect 2134 474 2203 507
rect 2634 474 2703 507
rect 3134 474 3203 507
rect 3634 474 3703 507
rect 4134 474 4203 507
rect 4634 474 4703 507
rect 5134 474 5203 507
<< obsli1 >>
rect 1012 4278 1212 4295
rect 1512 4278 1712 4295
rect 1218 4053 1235 4257
rect 1718 4053 1735 4257
rect 10720 4244 10789 4460
rect 1012 4014 1212 4031
rect 1512 4014 1712 4031
rect 1012 3908 1212 3925
rect 1512 3908 1712 3925
rect 1218 3683 1235 3887
rect 1718 3683 1735 3887
rect 1012 3644 1212 3661
rect 1512 3644 1712 3661
rect 5871 3448 6071 3465
rect 6321 3448 6521 3465
rect 6771 3448 6971 3465
rect 7221 3448 7421 3465
rect 7671 3448 7871 3465
rect 8121 3448 8321 3465
rect 8571 3448 8771 3465
rect 9021 3448 9221 3465
rect 5871 3184 6071 3201
rect 6321 3184 6521 3201
rect 6771 3184 6971 3201
rect 7221 3184 7421 3201
rect 7671 3184 7871 3201
rect 8121 3184 8321 3201
rect 8571 3184 8771 3201
rect 9021 3184 9221 3201
rect 5871 3078 6071 3095
rect 6321 3078 6521 3095
rect 6771 3078 6971 3095
rect 7221 3078 7421 3095
rect 7671 3078 7871 3095
rect 8121 3078 8321 3095
rect 8571 3078 8771 3095
rect 9021 3078 9221 3095
rect -2084 2938 -2015 2971
rect -1734 2938 -1665 2971
rect -1384 2938 -1315 2971
rect -1034 2938 -965 2971
rect -684 2938 -615 2971
rect -334 2938 -265 2971
rect 16 2938 85 2971
rect 366 2938 435 2971
rect 716 2938 785 2971
rect 1066 2938 1135 2971
rect 1916 2938 1985 2971
rect 2266 2938 2335 2971
rect 2616 2938 2685 2971
rect 2966 2938 3035 2971
rect 3316 2938 3385 2971
rect 3666 2938 3735 2971
rect 4016 2938 4085 2971
rect 4366 2938 4435 2971
rect 4716 2938 4785 2971
rect 5066 2938 5135 2971
rect -2127 1813 -2110 2817
rect -1998 1813 -1981 2817
rect -1777 1813 -1760 2817
rect -1648 1813 -1631 2817
rect -1427 1813 -1410 2817
rect -1298 1813 -1281 2817
rect -1077 1813 -1060 2817
rect -948 1813 -931 2817
rect -727 1813 -710 2817
rect -598 1813 -581 2817
rect -377 1813 -360 2817
rect -248 1813 -231 2817
rect -27 1813 -10 2817
rect 102 1813 119 2817
rect 323 1813 340 2817
rect 452 1813 469 2817
rect 673 1813 690 2817
rect 802 1813 819 2817
rect 1023 1813 1040 2817
rect 1152 1813 1169 2817
rect 1873 1813 1890 2817
rect 2002 1813 2019 2817
rect 2223 1813 2240 2817
rect 2352 1813 2369 2817
rect 2573 1813 2590 2817
rect 2702 1813 2719 2817
rect 2923 1813 2940 2817
rect 3052 1813 3069 2817
rect 3273 1813 3290 2817
rect 3402 1813 3419 2817
rect 3623 1813 3640 2817
rect 3752 1813 3769 2817
rect 3973 1813 3990 2817
rect 4102 1813 4119 2817
rect 4323 1813 4340 2817
rect 4452 1813 4469 2817
rect 4673 1813 4690 2817
rect 4802 1813 4819 2817
rect 5023 1813 5040 2817
rect 5152 1813 5169 2817
rect 5871 2814 6071 2831
rect 6321 2814 6521 2831
rect 6771 2814 6971 2831
rect 7221 2814 7421 2831
rect 7671 2814 7871 2831
rect 8121 2814 8321 2831
rect 8571 2814 8771 2831
rect 9021 2814 9221 2831
rect 1273 856 1290 960
rect 1273 606 1290 710
<< metal1 >>
rect -4600 4476 2133 4535
rect 920 4395 986 4476
rect 1420 4395 1486 4476
rect 920 4343 1150 4395
rect 1420 4343 1650 4395
rect 920 4255 986 4343
rect 920 4055 1009 4255
rect 920 3885 986 4055
rect 920 3685 1009 3885
rect 920 3592 986 3685
rect 920 3540 1150 3592
rect 1420 4255 1486 4343
rect 1420 4055 1509 4255
rect 1420 3885 1486 4055
rect 1420 3685 1509 3885
rect 1420 3592 1486 3685
rect 1420 3540 1650 3592
rect 2063 3737 2133 4476
rect 2063 3646 8995 3737
rect 5779 3565 5845 3646
rect 6229 3565 6295 3646
rect 6679 3565 6745 3646
rect 7129 3565 7195 3646
rect 7579 3565 7645 3646
rect 8029 3565 8095 3646
rect 8479 3565 8545 3646
rect 8929 3565 8995 3646
rect 5779 3513 6009 3565
rect 6229 3513 6459 3565
rect 6679 3513 6909 3565
rect 7129 3513 7359 3565
rect 7579 3513 7809 3565
rect 8029 3513 8259 3565
rect 8479 3513 8709 3565
rect 8929 3513 9159 3565
rect 5779 3425 5845 3513
rect 6097 3425 6164 3490
rect 5779 3225 5868 3425
rect 6074 3225 6164 3425
rect -2397 2971 -2345 2977
rect -2397 2945 -2384 2971
rect -2358 2945 -2345 2971
rect -2397 2939 -2345 2945
rect -2397 2913 -2384 2939
rect -2358 2913 -2345 2939
rect -2397 1376 -2345 2913
rect -2102 2831 -2006 2854
rect -1752 2831 -1656 2854
rect -1402 2831 -1306 2854
rect -1052 2831 -956 2854
rect -702 2831 -606 2854
rect -352 2831 -256 2854
rect -2 2831 94 2854
rect 348 2831 444 2854
rect 698 2831 794 2854
rect 1048 2831 1144 2854
rect 1898 2831 1994 2854
rect 2248 2831 2344 2854
rect 2598 2831 2694 2854
rect 2948 2831 3044 2854
rect 3298 2831 3394 2854
rect 3648 2831 3744 2854
rect 3998 2831 4094 2854
rect 4348 2831 4444 2854
rect 4698 2831 4794 2854
rect 5779 3055 5845 3225
rect 6097 3055 6164 3225
rect 5779 2855 5868 3055
rect 6074 2855 6164 3055
rect 5048 2831 5144 2854
rect 5779 2762 5845 2855
rect 5779 2710 6009 2762
rect 6097 2625 6164 2855
rect 6229 3425 6295 3513
rect 6547 3425 6614 3490
rect 6229 3225 6318 3425
rect 6524 3225 6614 3425
rect 6229 3055 6295 3225
rect 6547 3055 6614 3225
rect 6229 2855 6318 3055
rect 6524 2855 6614 3055
rect 6229 2762 6295 2855
rect 6229 2710 6459 2762
rect 6547 2625 6614 2855
rect 6679 3425 6745 3513
rect 6997 3425 7064 3490
rect 6679 3225 6768 3425
rect 6974 3225 7064 3425
rect 6679 3055 6745 3225
rect 6997 3055 7064 3225
rect 6679 2855 6768 3055
rect 6974 2855 7064 3055
rect 6679 2762 6745 2855
rect 6679 2710 6909 2762
rect 6997 2625 7064 2855
rect 7129 3425 7195 3513
rect 7447 3425 7514 3490
rect 7129 3225 7218 3425
rect 7424 3225 7514 3425
rect 7129 3055 7195 3225
rect 7447 3055 7514 3225
rect 7129 2855 7218 3055
rect 7424 2855 7514 3055
rect 7129 2762 7195 2855
rect 7129 2710 7359 2762
rect 7447 2625 7514 2855
rect 7579 3425 7645 3513
rect 7897 3425 7964 3490
rect 7579 3225 7668 3425
rect 7874 3225 7964 3425
rect 7579 3055 7645 3225
rect 7897 3055 7964 3225
rect 7579 2855 7668 3055
rect 7874 2855 7964 3055
rect 7579 2762 7645 2855
rect 7579 2710 7809 2762
rect 7897 2625 7964 2855
rect 8029 3425 8095 3513
rect 8347 3425 8414 3490
rect 8029 3225 8118 3425
rect 8324 3225 8414 3425
rect 8029 3055 8095 3225
rect 8347 3055 8414 3225
rect 8029 2855 8118 3055
rect 8324 2855 8414 3055
rect 8029 2762 8095 2855
rect 8029 2710 8259 2762
rect 8347 2625 8414 2855
rect 8479 3425 8545 3513
rect 8797 3425 8864 3490
rect 8479 3225 8568 3425
rect 8774 3225 8864 3425
rect 8479 3055 8545 3225
rect 8797 3055 8864 3225
rect 8479 2855 8568 3055
rect 8774 2855 8864 3055
rect 8479 2762 8545 2855
rect 8479 2710 8709 2762
rect 8797 2625 8864 2855
rect 8929 3425 8995 3513
rect 9247 3425 9314 3490
rect 8929 3225 9018 3425
rect 9224 3225 9314 3425
rect 8929 3055 8995 3225
rect 9247 3055 9314 3225
rect 8929 2855 9018 3055
rect 9224 2855 9314 3055
rect 10537 2991 10578 3814
rect 10537 2965 10545 2991
rect 10571 2965 10578 2991
rect 10537 2959 10578 2965
rect 10537 2933 10545 2959
rect 10571 2933 10578 2959
rect 10537 2927 10578 2933
rect 8929 2762 8995 2855
rect 8929 2710 9159 2762
rect 9247 2625 9314 2855
rect 6097 2532 9314 2625
rect -2102 1742 -2006 1799
rect -2102 1716 -2083 1742
rect -2057 1716 -2051 1742
rect -2025 1716 -2006 1742
rect -2102 1679 -2006 1716
rect -1752 1742 -1656 1799
rect -1752 1716 -1733 1742
rect -1707 1716 -1701 1742
rect -1675 1716 -1656 1742
rect -1752 1679 -1656 1716
rect -1402 1742 -1306 1799
rect -1402 1716 -1383 1742
rect -1357 1716 -1351 1742
rect -1325 1716 -1306 1742
rect -1402 1679 -1306 1716
rect -1052 1742 -956 1799
rect -1052 1716 -1033 1742
rect -1007 1716 -1001 1742
rect -975 1716 -956 1742
rect -1052 1679 -956 1716
rect -702 1742 -606 1799
rect -702 1716 -683 1742
rect -657 1716 -651 1742
rect -625 1716 -606 1742
rect -702 1679 -606 1716
rect -352 1742 -256 1799
rect -352 1716 -333 1742
rect -307 1716 -301 1742
rect -275 1716 -256 1742
rect -352 1679 -256 1716
rect -2 1742 94 1799
rect -2 1716 18 1742
rect 44 1716 50 1742
rect 76 1716 94 1742
rect -2 1679 94 1716
rect 348 1742 444 1799
rect 348 1716 368 1742
rect 394 1716 400 1742
rect 426 1716 444 1742
rect 348 1679 444 1716
rect 698 1742 794 1799
rect 698 1716 718 1742
rect 744 1716 750 1742
rect 776 1716 794 1742
rect 698 1679 794 1716
rect 1048 1742 1144 1799
rect 1048 1716 1068 1742
rect 1094 1716 1100 1742
rect 1126 1716 1144 1742
rect 1048 1679 1144 1716
rect 1898 1742 1994 1799
rect 1898 1716 1918 1742
rect 1944 1716 1950 1742
rect 1976 1716 1994 1742
rect 1898 1679 1994 1716
rect 2248 1742 2344 1799
rect 2248 1716 2268 1742
rect 2294 1716 2300 1742
rect 2326 1716 2344 1742
rect 2248 1679 2344 1716
rect 2598 1742 2694 1799
rect 2598 1716 2618 1742
rect 2644 1716 2650 1742
rect 2676 1716 2694 1742
rect 2598 1679 2694 1716
rect 2948 1742 3044 1799
rect 2948 1716 2968 1742
rect 2994 1716 3000 1742
rect 3026 1716 3044 1742
rect 2948 1679 3044 1716
rect 3298 1742 3394 1799
rect 3298 1716 3318 1742
rect 3344 1716 3350 1742
rect 3376 1716 3394 1742
rect 3298 1679 3394 1716
rect 3648 1742 3744 1799
rect 3648 1716 3668 1742
rect 3694 1716 3700 1742
rect 3726 1716 3744 1742
rect 3648 1679 3744 1716
rect 3998 1742 4094 1799
rect 3998 1716 4018 1742
rect 4044 1716 4050 1742
rect 4076 1716 4094 1742
rect 3998 1679 4094 1716
rect 4348 1742 4444 1799
rect 4348 1716 4368 1742
rect 4394 1716 4400 1742
rect 4426 1716 4444 1742
rect 4348 1679 4444 1716
rect 4698 1742 4794 1799
rect 4698 1716 4718 1742
rect 4744 1716 4750 1742
rect 4776 1716 4794 1742
rect 4698 1679 4794 1716
rect 5048 1742 5144 1799
rect 5048 1716 5068 1742
rect 5094 1716 5100 1742
rect 5126 1716 5144 1742
rect 5048 1679 5144 1716
rect 6146 1988 6231 2532
rect 10725 1988 10784 3242
rect 6146 1870 16925 1988
rect -2397 1350 -2384 1376
rect -2358 1350 -2345 1376
rect -2397 1344 -2345 1350
rect -2397 1318 -2384 1344
rect -2358 1318 -2345 1344
rect -2397 1307 -2345 1318
rect -4600 1144 856 1206
rect 637 1071 702 1073
rect 479 1044 702 1071
rect 479 1038 701 1044
rect 479 958 541 1038
rect 569 974 765 997
rect 793 958 856 1144
rect 1137 1071 1202 1073
rect 479 858 564 958
rect 770 858 856 958
rect 479 708 541 858
rect 569 819 765 842
rect 793 819 856 858
rect 569 797 856 819
rect 569 771 642 797
rect 668 771 674 797
rect 700 771 856 797
rect 569 747 856 771
rect 569 724 765 747
rect 793 708 856 747
rect 479 608 564 708
rect 770 608 856 708
rect 479 505 541 608
rect 569 569 765 592
rect 479 472 701 505
rect 479 357 541 472
rect 793 430 856 608
rect 979 1044 1202 1071
rect 979 1038 1201 1044
rect 979 958 1041 1038
rect 1069 974 1265 997
rect 6146 1260 6231 1870
rect 1793 1199 6231 1260
rect 1637 1071 1702 1073
rect 979 858 1064 958
rect 979 708 1041 858
rect 1069 797 1265 842
rect 1069 771 1142 797
rect 1168 771 1174 797
rect 1200 771 1265 797
rect 1069 724 1265 771
rect 979 608 1064 708
rect 979 505 1041 608
rect 1069 569 1265 592
rect 979 472 1201 505
rect 979 357 1041 472
rect 1479 1044 1702 1071
rect 1479 1038 1701 1044
rect 1479 958 1541 1038
rect 1569 974 1765 997
rect 1793 958 1856 1199
rect 2137 1071 2202 1073
rect 1479 858 1564 958
rect 1770 858 1856 958
rect 1479 708 1541 858
rect 1569 797 1765 842
rect 1569 771 1642 797
rect 1668 771 1674 797
rect 1700 771 1765 797
rect 1569 724 1765 771
rect 1793 708 1856 858
rect 1479 608 1564 708
rect 1770 608 1856 708
rect 1479 505 1541 608
rect 1569 569 1765 592
rect 1479 472 1701 505
rect 1479 357 1541 472
rect 1793 430 1856 608
rect 1979 1044 2202 1071
rect 1979 1038 2201 1044
rect 1979 958 2041 1038
rect 2069 974 2265 997
rect 2293 958 2356 1199
rect 2637 1071 2702 1073
rect 1979 858 2064 958
rect 2270 858 2356 958
rect 1979 708 2041 858
rect 2069 797 2265 842
rect 2069 771 2142 797
rect 2168 771 2174 797
rect 2200 771 2265 797
rect 2069 724 2265 771
rect 2293 708 2356 858
rect 1979 608 2064 708
rect 2270 608 2356 708
rect 1979 505 2041 608
rect 2069 569 2265 592
rect 1979 472 2201 505
rect 1979 357 2041 472
rect 2293 430 2356 608
rect 2479 1044 2702 1071
rect 2479 1038 2701 1044
rect 2479 958 2541 1038
rect 2569 974 2765 997
rect 2793 958 2856 1199
rect 3137 1071 3202 1073
rect 2479 858 2564 958
rect 2770 858 2856 958
rect 2479 708 2541 858
rect 2569 797 2765 842
rect 2569 771 2642 797
rect 2668 771 2674 797
rect 2700 771 2765 797
rect 2569 724 2765 771
rect 2793 708 2856 858
rect 2479 608 2564 708
rect 2770 608 2856 708
rect 2479 505 2541 608
rect 2569 569 2765 592
rect 2479 472 2701 505
rect 2479 357 2541 472
rect 2793 430 2856 608
rect 2979 1044 3202 1071
rect 2979 1038 3201 1044
rect 2979 958 3041 1038
rect 3069 974 3265 997
rect 3293 958 3356 1199
rect 3637 1071 3702 1073
rect 2979 858 3064 958
rect 3270 858 3356 958
rect 2979 708 3041 858
rect 3069 797 3265 842
rect 3069 771 3142 797
rect 3168 771 3174 797
rect 3200 771 3265 797
rect 3069 724 3265 771
rect 3293 708 3356 858
rect 2979 608 3064 708
rect 3270 608 3356 708
rect 2979 505 3041 608
rect 3069 569 3265 592
rect 2979 472 3201 505
rect 2979 357 3041 472
rect 3293 430 3356 608
rect 3479 1044 3702 1071
rect 3479 1038 3701 1044
rect 3479 958 3541 1038
rect 3569 974 3765 997
rect 3793 958 3856 1199
rect 4137 1071 4202 1073
rect 3479 858 3564 958
rect 3770 858 3856 958
rect 3479 708 3541 858
rect 3569 797 3765 842
rect 3569 771 3642 797
rect 3668 771 3674 797
rect 3700 771 3765 797
rect 3569 724 3765 771
rect 3793 708 3856 858
rect 3479 608 3564 708
rect 3770 608 3856 708
rect 3479 505 3541 608
rect 3569 569 3765 592
rect 3479 472 3701 505
rect 3479 357 3541 472
rect 3793 430 3856 608
rect 3979 1044 4202 1071
rect 3979 1038 4201 1044
rect 3979 958 4041 1038
rect 4069 974 4265 997
rect 4293 958 4356 1199
rect 4637 1071 4702 1073
rect 3979 858 4064 958
rect 4270 858 4356 958
rect 3979 708 4041 858
rect 4069 797 4265 842
rect 4069 771 4142 797
rect 4168 771 4174 797
rect 4200 771 4265 797
rect 4069 724 4265 771
rect 4293 708 4356 858
rect 3979 608 4064 708
rect 4270 608 4356 708
rect 3979 505 4041 608
rect 4069 569 4265 592
rect 3979 472 4201 505
rect 3979 357 4041 472
rect 4293 430 4356 608
rect 4479 1044 4702 1071
rect 4479 1038 4701 1044
rect 4479 958 4541 1038
rect 4569 974 4765 997
rect 4793 958 4856 1199
rect 5137 1071 5202 1073
rect 4479 858 4564 958
rect 4770 858 4856 958
rect 4479 708 4541 858
rect 4569 797 4765 842
rect 4569 771 4642 797
rect 4668 771 4674 797
rect 4700 771 4765 797
rect 4569 724 4765 771
rect 4793 708 4856 858
rect 4479 608 4564 708
rect 4770 608 4856 708
rect 4479 505 4541 608
rect 4569 569 4765 592
rect 4479 472 4701 505
rect 4479 357 4541 472
rect 4793 430 4856 608
rect 4979 1044 5202 1071
rect 4979 1038 5201 1044
rect 4979 958 5041 1038
rect 5069 974 5265 997
rect 5293 958 5356 1199
rect 4979 858 5064 958
rect 5270 858 5356 958
rect 4979 708 5041 858
rect 5069 797 5265 842
rect 5069 771 5142 797
rect 5168 771 5174 797
rect 5200 771 5265 797
rect 5069 724 5265 771
rect 5293 708 5356 858
rect 4979 608 5064 708
rect 5270 608 5356 708
rect 4979 505 5041 608
rect 5069 569 5265 592
rect 4979 472 5201 505
rect 4979 357 5041 472
rect 5293 430 5356 608
rect -4600 332 5409 357
rect -4600 306 -2384 332
rect -2358 306 5409 332
rect -4600 300 5409 306
rect -4600 274 -2384 300
rect -2358 274 5409 300
rect -4600 248 5409 274
<< via1 >>
rect -2384 2945 -2358 2971
rect -2384 2913 -2358 2939
rect 10545 2965 10571 2991
rect 10545 2933 10571 2959
rect -2083 1716 -2057 1742
rect -2051 1716 -2025 1742
rect -1733 1716 -1707 1742
rect -1701 1716 -1675 1742
rect -1383 1716 -1357 1742
rect -1351 1716 -1325 1742
rect -1033 1716 -1007 1742
rect -1001 1716 -975 1742
rect -683 1716 -657 1742
rect -651 1716 -625 1742
rect -333 1716 -307 1742
rect -301 1716 -275 1742
rect 18 1716 44 1742
rect 50 1716 76 1742
rect 368 1716 394 1742
rect 400 1716 426 1742
rect 718 1716 744 1742
rect 750 1716 776 1742
rect 1068 1716 1094 1742
rect 1100 1716 1126 1742
rect 1918 1716 1944 1742
rect 1950 1716 1976 1742
rect 2268 1716 2294 1742
rect 2300 1716 2326 1742
rect 2618 1716 2644 1742
rect 2650 1716 2676 1742
rect 2968 1716 2994 1742
rect 3000 1716 3026 1742
rect 3318 1716 3344 1742
rect 3350 1716 3376 1742
rect 3668 1716 3694 1742
rect 3700 1716 3726 1742
rect 4018 1716 4044 1742
rect 4050 1716 4076 1742
rect 4368 1716 4394 1742
rect 4400 1716 4426 1742
rect 4718 1716 4744 1742
rect 4750 1716 4776 1742
rect 5068 1716 5094 1742
rect 5100 1716 5126 1742
rect -2384 1350 -2358 1376
rect -2384 1318 -2358 1344
rect 642 771 668 797
rect 674 771 700 797
rect 1142 771 1168 797
rect 1174 771 1200 797
rect 1642 771 1668 797
rect 1674 771 1700 797
rect 2142 771 2168 797
rect 2174 771 2200 797
rect 2642 771 2668 797
rect 2674 771 2700 797
rect 3142 771 3168 797
rect 3174 771 3200 797
rect 3642 771 3668 797
rect 3674 771 3700 797
rect 4142 771 4168 797
rect 4174 771 4200 797
rect 4642 771 4668 797
rect 4674 771 4700 797
rect 5142 771 5168 797
rect 5174 771 5200 797
rect -2384 306 -2358 332
rect -2384 274 -2358 300
<< obsm1 >>
rect 1014 4275 1210 4298
rect 1238 4255 1305 4320
rect 1215 4055 1305 4255
rect 1014 4011 1210 4034
rect 1238 4011 1305 4055
rect 1014 3928 1305 4011
rect 1014 3905 1210 3928
rect 1238 3885 1305 3928
rect 1215 3685 1305 3885
rect 1014 3641 1210 3664
rect 1238 3207 1305 3685
rect 1514 4275 1710 4298
rect 1738 4255 1805 4320
rect 1715 4055 1805 4255
rect 1514 3905 1710 4034
rect 1738 3885 1805 4055
rect 1715 3685 1805 3885
rect 1514 3641 1710 3664
rect 1006 3170 1307 3207
rect 1738 3205 1805 3685
rect 10725 4247 10784 4457
rect -2198 3091 1307 3170
rect 1739 3170 1805 3205
rect 5873 3445 6069 3468
rect 1739 3155 5020 3170
rect 1739 3123 5030 3155
rect 1739 3094 5020 3123
rect -2198 3090 1020 3091
rect -2198 2815 -2130 3090
rect -1848 2815 -1780 3090
rect -1498 2815 -1430 3090
rect -1148 2815 -1080 3090
rect -798 2815 -730 3090
rect -448 2815 -380 3090
rect -98 2815 -30 3090
rect 252 2815 320 3090
rect 602 2815 670 3090
rect 952 2815 1020 3090
rect 1802 3090 5020 3094
rect 1802 2815 1870 3090
rect 2152 2815 2220 3090
rect 2502 2815 2570 3090
rect 2852 2815 2920 3090
rect 3202 2815 3270 3090
rect 3552 2815 3620 3090
rect 3902 2815 3970 3090
rect 4252 2815 4320 3090
rect 4602 2815 4670 3090
rect 4952 2815 5020 3090
rect 5873 3075 6069 3204
rect -2198 1815 -2107 2815
rect -2001 1815 -1910 2815
rect -1848 1815 -1757 2815
rect -1651 1815 -1560 2815
rect -1498 1815 -1407 2815
rect -1301 1815 -1210 2815
rect -1148 1815 -1057 2815
rect -951 1815 -860 2815
rect -798 1815 -707 2815
rect -601 1815 -510 2815
rect -448 1815 -357 2815
rect -251 1815 -160 2815
rect -98 1815 -7 2815
rect 99 1815 190 2815
rect 252 1815 343 2815
rect 449 1815 540 2815
rect 602 1815 693 2815
rect 799 1815 890 2815
rect 952 1815 1043 2815
rect 1149 1815 1240 2815
rect 1802 1815 1893 2815
rect 1999 1815 2090 2815
rect 2152 1815 2243 2815
rect 2349 1815 2440 2815
rect 2502 1815 2593 2815
rect 2699 1815 2790 2815
rect 2852 1815 2943 2815
rect 3049 1815 3140 2815
rect 3202 1815 3293 2815
rect 3399 1815 3490 2815
rect 3552 1815 3643 2815
rect 3749 1815 3840 2815
rect 3902 1815 3993 2815
rect 4099 1815 4190 2815
rect 4252 1815 4343 2815
rect 4449 1815 4540 2815
rect 4602 1815 4693 2815
rect 4799 1815 4890 2815
rect 4952 1815 5043 2815
rect 5149 1815 5240 2815
rect 5873 2811 6069 2834
rect 6323 3445 6519 3468
rect 6323 3075 6519 3204
rect 6323 2811 6519 2834
rect 6773 3445 6969 3468
rect 6773 3075 6969 3204
rect 6773 2811 6969 2834
rect 7223 3445 7419 3468
rect 7223 3075 7419 3204
rect 7223 2811 7419 2834
rect 7673 3445 7869 3468
rect 7673 3075 7869 3204
rect 7673 2811 7869 2834
rect 8123 3445 8319 3468
rect 8123 3075 8319 3204
rect 8123 2811 8319 2834
rect 8573 3445 8769 3468
rect 8573 3075 8769 3204
rect 8573 2811 8769 2834
rect 9023 3445 9219 3468
rect 9023 3075 9219 3204
rect 9023 2811 9219 2834
rect -1978 1540 -1910 1815
rect -1628 1540 -1560 1815
rect -1278 1540 -1210 1815
rect -928 1540 -860 1815
rect -578 1540 -510 1815
rect -228 1540 -160 1815
rect 122 1540 190 1815
rect 472 1540 540 1815
rect 822 1540 890 1815
rect 1172 1540 1240 1815
rect 2022 1540 2090 1815
rect 2372 1540 2440 1815
rect 2722 1540 2790 1815
rect 3072 1540 3140 1815
rect 3422 1540 3490 1815
rect 3772 1540 3840 1815
rect 4122 1540 4190 1815
rect 4472 1540 4540 1815
rect 4822 1540 4890 1815
rect 5172 1540 5240 1815
rect -1978 1460 5240 1540
rect 1293 958 1356 1460
rect 1270 858 1356 958
rect 1293 708 1356 858
rect 1270 608 1356 708
rect 1293 430 1356 608
<< metal2 >>
rect 10542 2991 10574 2994
rect 10542 2977 10545 2991
rect -2397 2971 10545 2977
rect -2397 2945 -2384 2971
rect -2358 2965 10545 2971
rect 10571 2977 10574 2991
rect 10571 2965 10578 2977
rect -2358 2959 10578 2965
rect -2358 2945 10545 2959
rect -2397 2939 10545 2945
rect -2397 2927 -2384 2939
rect -2387 2913 -2384 2927
rect -2358 2933 10545 2939
rect 10571 2933 10578 2959
rect -2358 2927 10578 2933
rect -2358 2913 -2355 2927
rect -2387 2910 -2355 2913
rect -4600 1742 1137 1750
rect -4600 1716 -2083 1742
rect -2057 1716 -2051 1742
rect -2025 1716 -1733 1742
rect -1707 1716 -1701 1742
rect -1675 1716 -1383 1742
rect -1357 1716 -1351 1742
rect -1325 1716 -1033 1742
rect -1007 1716 -1001 1742
rect -975 1716 -683 1742
rect -657 1716 -651 1742
rect -625 1716 -333 1742
rect -307 1716 -301 1742
rect -275 1716 18 1742
rect 44 1716 50 1742
rect 76 1716 368 1742
rect 394 1716 400 1742
rect 426 1716 718 1742
rect 744 1716 750 1742
rect 776 1716 1068 1742
rect 1094 1716 1100 1742
rect 1126 1716 1137 1742
rect -4600 1707 1137 1716
rect 1910 1742 16925 1750
rect 1910 1716 1918 1742
rect 1944 1716 1950 1742
rect 1976 1716 2268 1742
rect 2294 1716 2300 1742
rect 2326 1716 2618 1742
rect 2644 1716 2650 1742
rect 2676 1716 2968 1742
rect 2994 1716 3000 1742
rect 3026 1716 3318 1742
rect 3344 1716 3350 1742
rect 3376 1716 3668 1742
rect 3694 1716 3700 1742
rect 3726 1716 4018 1742
rect 4044 1716 4050 1742
rect 4076 1716 4368 1742
rect 4394 1716 4400 1742
rect 4426 1716 4718 1742
rect 4744 1716 4750 1742
rect 4776 1716 5068 1742
rect 5094 1716 5100 1742
rect 5126 1716 16925 1742
rect 1910 1707 16925 1716
rect -2390 1376 -2351 1381
rect -2390 1350 -2384 1376
rect -2358 1350 -2351 1376
rect -2390 1344 -2351 1350
rect -2390 1318 -2384 1344
rect -2358 1318 -2351 1344
rect -2390 332 -2351 1318
rect 634 797 5214 805
rect 634 771 642 797
rect 668 771 674 797
rect 700 771 1142 797
rect 1168 771 1174 797
rect 1200 771 1642 797
rect 1668 771 1674 797
rect 1700 771 2142 797
rect 2168 771 2174 797
rect 2200 771 2642 797
rect 2668 771 2674 797
rect 2700 771 3142 797
rect 3168 771 3174 797
rect 3200 771 3642 797
rect 3668 771 3674 797
rect 3700 771 4142 797
rect 4168 771 4174 797
rect 4200 771 4642 797
rect 4668 771 4674 797
rect 4700 771 5142 797
rect 5168 771 5174 797
rect 5200 771 5214 797
rect 634 763 5214 771
rect -2390 306 -2384 332
rect -2358 306 -2351 332
rect -2390 300 -2351 306
rect -2390 274 -2384 300
rect -2358 274 -2351 300
rect -2390 254 -2351 274
<< obsm2 >>
rect 1082 3952 1652 3990
rect 5837 3165 5919 8561
rect 10730 4372 10778 4453
rect 4940 3115 9166 3165
<< obsm3 >>
rect 5859 8554 5897 8556
rect 5854 8463 5902 8554
rect -4360 5185 -1260 8334
rect -860 5185 2241 8334
rect 2641 5185 5741 8334
rect 6141 5185 9241 8334
rect 9641 5185 12741 8334
rect 13141 5185 16241 8334
rect 10735 4454 10773 4458
rect 10729 4370 10779 4454
rect 10735 4365 10773 4370
<< obsm4 >>
rect -4290 8437 16171 8609
rect -4290 5304 -1329 8265
rect -790 5304 2171 8265
rect 2710 5304 5671 8265
rect 6210 5304 9171 8265
rect 9710 5304 12671 8265
rect 13210 5304 16171 8265
rect -4354 5187 -1266 5235
rect -854 5187 2235 5235
rect 2647 5187 5735 5235
rect 6147 5187 9235 5235
rect 9647 5187 12735 5235
rect 13147 5187 16235 5235
rect -4354 5091 16235 5187
rect 10735 4365 10773 5091
<< obsm5 >>
rect -4149 8077 -3847 8594
rect -649 8077 -347 8594
rect 2851 8077 3153 8594
rect 6351 8077 6653 8594
rect 9851 8077 10153 8594
rect 13351 8077 13653 8594
<< labels >>
rlabel metal2 s -2390 254 -2351 1381 4 vss
port 1 nsew
rlabel metal2 s -2387 2910 -2355 2927 4 vss
port 1 nsew
rlabel metal2 s -2397 2927 10578 2977 6 vss
port 1 nsew
rlabel metal2 s 10542 2977 10574 2994 6 vss
port 1 nsew
rlabel via1 s -2384 274 -2358 300 4 vss
port 1 nsew
rlabel via1 s -2384 306 -2358 332 4 vss
port 1 nsew
rlabel via1 s -2384 1318 -2358 1344 4 vss
port 1 nsew
rlabel via1 s -2384 1350 -2358 1376 4 vss
port 1 nsew
rlabel via1 s 10545 2933 10571 2959 6 vss
port 1 nsew
rlabel via1 s 10545 2965 10571 2991 6 vss
port 1 nsew
rlabel via1 s -2384 2913 -2358 2939 4 vss
port 1 nsew
rlabel via1 s -2384 2945 -2358 2971 4 vss
port 1 nsew
rlabel metal1 s -4600 248 5409 357 6 vss
port 1 nsew
rlabel metal1 s 4979 357 5041 472 6 vss
port 1 nsew
rlabel metal1 s 4479 357 4541 472 6 vss
port 1 nsew
rlabel metal1 s 3979 357 4041 472 6 vss
port 1 nsew
rlabel metal1 s 3479 357 3541 472 6 vss
port 1 nsew
rlabel metal1 s 2979 357 3041 472 6 vss
port 1 nsew
rlabel metal1 s 2479 357 2541 472 6 vss
port 1 nsew
rlabel metal1 s 1979 357 2041 472 6 vss
port 1 nsew
rlabel metal1 s 1479 357 1541 472 6 vss
port 1 nsew
rlabel metal1 s 979 357 1041 472 6 vss
port 1 nsew
rlabel metal1 s 479 357 541 472 6 vss
port 1 nsew
rlabel metal1 s 4979 472 5201 476 6 vss
port 1 nsew
rlabel metal1 s 4479 472 4701 476 6 vss
port 1 nsew
rlabel metal1 s 3979 472 4201 476 6 vss
port 1 nsew
rlabel metal1 s 3479 472 3701 476 6 vss
port 1 nsew
rlabel metal1 s 2979 472 3201 476 6 vss
port 1 nsew
rlabel metal1 s 2479 472 2701 476 6 vss
port 1 nsew
rlabel metal1 s 1979 472 2201 476 6 vss
port 1 nsew
rlabel metal1 s 1479 472 1701 476 6 vss
port 1 nsew
rlabel metal1 s 979 472 1201 476 6 vss
port 1 nsew
rlabel metal1 s 479 472 701 476 6 vss
port 1 nsew
rlabel metal1 s 4979 476 5201 505 6 vss
port 1 nsew
rlabel metal1 s 4479 476 4701 505 6 vss
port 1 nsew
rlabel metal1 s 3979 476 4201 505 6 vss
port 1 nsew
rlabel metal1 s 3479 476 3701 505 6 vss
port 1 nsew
rlabel metal1 s 2979 476 3201 505 6 vss
port 1 nsew
rlabel metal1 s 2479 476 2701 505 6 vss
port 1 nsew
rlabel metal1 s 1979 476 2201 505 6 vss
port 1 nsew
rlabel metal1 s 1479 476 1701 505 6 vss
port 1 nsew
rlabel metal1 s 979 476 1201 505 6 vss
port 1 nsew
rlabel metal1 s 479 476 701 505 6 vss
port 1 nsew
rlabel metal1 s 4979 505 5201 505 6 vss
port 1 nsew
rlabel metal1 s 4479 505 4701 505 6 vss
port 1 nsew
rlabel metal1 s 3979 505 4201 505 6 vss
port 1 nsew
rlabel metal1 s 3479 505 3701 505 6 vss
port 1 nsew
rlabel metal1 s 2979 505 3201 505 6 vss
port 1 nsew
rlabel metal1 s 2479 505 2701 505 6 vss
port 1 nsew
rlabel metal1 s 1979 505 2201 505 6 vss
port 1 nsew
rlabel metal1 s 1479 505 1701 505 6 vss
port 1 nsew
rlabel metal1 s 979 505 1201 505 6 vss
port 1 nsew
rlabel metal1 s 479 505 701 505 6 vss
port 1 nsew
rlabel metal1 s 4979 505 5041 608 6 vss
port 1 nsew
rlabel metal1 s 4479 505 4541 608 6 vss
port 1 nsew
rlabel metal1 s 3979 505 4041 608 6 vss
port 1 nsew
rlabel metal1 s 3479 505 3541 608 6 vss
port 1 nsew
rlabel metal1 s 2979 505 3041 608 6 vss
port 1 nsew
rlabel metal1 s 2479 505 2541 608 6 vss
port 1 nsew
rlabel metal1 s 1979 505 2041 608 6 vss
port 1 nsew
rlabel metal1 s 1479 505 1541 608 6 vss
port 1 nsew
rlabel metal1 s 979 505 1041 608 6 vss
port 1 nsew
rlabel metal1 s 479 505 541 608 6 vss
port 1 nsew
rlabel metal1 s 4979 608 5064 708 6 vss
port 1 nsew
rlabel metal1 s 4479 608 4564 708 6 vss
port 1 nsew
rlabel metal1 s 3979 608 4064 708 6 vss
port 1 nsew
rlabel metal1 s 3479 608 3564 708 6 vss
port 1 nsew
rlabel metal1 s 2979 608 3064 708 6 vss
port 1 nsew
rlabel metal1 s 2479 608 2564 708 6 vss
port 1 nsew
rlabel metal1 s 1979 608 2064 708 6 vss
port 1 nsew
rlabel metal1 s 1479 608 1564 708 6 vss
port 1 nsew
rlabel metal1 s 979 608 1064 708 6 vss
port 1 nsew
rlabel metal1 s 479 608 564 708 6 vss
port 1 nsew
rlabel metal1 s 4979 708 5041 858 6 vss
port 1 nsew
rlabel metal1 s 4479 708 4541 858 6 vss
port 1 nsew
rlabel metal1 s 3979 708 4041 858 6 vss
port 1 nsew
rlabel metal1 s 3479 708 3541 858 6 vss
port 1 nsew
rlabel metal1 s 2979 708 3041 858 6 vss
port 1 nsew
rlabel metal1 s 2479 708 2541 858 6 vss
port 1 nsew
rlabel metal1 s 1979 708 2041 858 6 vss
port 1 nsew
rlabel metal1 s 1479 708 1541 858 6 vss
port 1 nsew
rlabel metal1 s 979 708 1041 858 6 vss
port 1 nsew
rlabel metal1 s 479 708 541 858 6 vss
port 1 nsew
rlabel metal1 s 4979 858 5064 958 6 vss
port 1 nsew
rlabel metal1 s 4479 858 4564 958 6 vss
port 1 nsew
rlabel metal1 s 3979 858 4064 958 6 vss
port 1 nsew
rlabel metal1 s 3479 858 3564 958 6 vss
port 1 nsew
rlabel metal1 s 2979 858 3064 958 6 vss
port 1 nsew
rlabel metal1 s 2479 858 2564 958 6 vss
port 1 nsew
rlabel metal1 s 1979 858 2064 958 6 vss
port 1 nsew
rlabel metal1 s 1479 858 1564 958 6 vss
port 1 nsew
rlabel metal1 s 979 858 1064 958 6 vss
port 1 nsew
rlabel metal1 s 479 858 564 958 6 vss
port 1 nsew
rlabel metal1 s 4979 958 5041 1038 6 vss
port 1 nsew
rlabel metal1 s 4479 958 4541 1038 6 vss
port 1 nsew
rlabel metal1 s 3979 958 4041 1038 6 vss
port 1 nsew
rlabel metal1 s 3479 958 3541 1038 6 vss
port 1 nsew
rlabel metal1 s 2979 958 3041 1038 6 vss
port 1 nsew
rlabel metal1 s 2479 958 2541 1038 6 vss
port 1 nsew
rlabel metal1 s 1979 958 2041 1038 6 vss
port 1 nsew
rlabel metal1 s 1479 958 1541 1038 6 vss
port 1 nsew
rlabel metal1 s 979 958 1041 1038 6 vss
port 1 nsew
rlabel metal1 s 479 958 541 1038 6 vss
port 1 nsew
rlabel metal1 s 4979 1038 5201 1044 6 vss
port 1 nsew
rlabel metal1 s 4479 1038 4701 1044 6 vss
port 1 nsew
rlabel metal1 s 3979 1038 4201 1044 6 vss
port 1 nsew
rlabel metal1 s 3479 1038 3701 1044 6 vss
port 1 nsew
rlabel metal1 s 2979 1038 3201 1044 6 vss
port 1 nsew
rlabel metal1 s 2479 1038 2701 1044 6 vss
port 1 nsew
rlabel metal1 s 1979 1038 2201 1044 6 vss
port 1 nsew
rlabel metal1 s 1479 1038 1701 1044 6 vss
port 1 nsew
rlabel metal1 s 979 1038 1201 1044 6 vss
port 1 nsew
rlabel metal1 s 479 1038 701 1044 6 vss
port 1 nsew
rlabel metal1 s 4979 1044 5202 1071 6 vss
port 1 nsew
rlabel metal1 s 4479 1044 4702 1071 6 vss
port 1 nsew
rlabel metal1 s 3979 1044 4202 1071 6 vss
port 1 nsew
rlabel metal1 s 3479 1044 3702 1071 6 vss
port 1 nsew
rlabel metal1 s 2979 1044 3202 1071 6 vss
port 1 nsew
rlabel metal1 s 2479 1044 2702 1071 6 vss
port 1 nsew
rlabel metal1 s 1979 1044 2202 1071 6 vss
port 1 nsew
rlabel metal1 s 1479 1044 1702 1071 6 vss
port 1 nsew
rlabel metal1 s 979 1044 1202 1071 6 vss
port 1 nsew
rlabel metal1 s 479 1044 702 1071 6 vss
port 1 nsew
rlabel metal1 s 5137 1071 5202 1073 6 vss
port 1 nsew
rlabel metal1 s 4637 1071 4702 1073 6 vss
port 1 nsew
rlabel metal1 s 4137 1071 4202 1073 6 vss
port 1 nsew
rlabel metal1 s 3637 1071 3702 1073 6 vss
port 1 nsew
rlabel metal1 s 3137 1071 3202 1073 6 vss
port 1 nsew
rlabel metal1 s 2637 1071 2702 1073 6 vss
port 1 nsew
rlabel metal1 s 2137 1071 2202 1073 6 vss
port 1 nsew
rlabel metal1 s 1637 1071 1702 1073 6 vss
port 1 nsew
rlabel metal1 s 1137 1071 1202 1073 6 vss
port 1 nsew
rlabel metal1 s 637 1071 702 1073 6 vss
port 1 nsew
rlabel metal1 s 10537 2927 10578 3814 6 vss
port 1 nsew
rlabel metal1 s -2397 1307 -2345 2977 4 vss
port 1 nsew
rlabel locali s 5134 474 5203 507 6 vss
port 1 nsew
rlabel locali s 4634 474 4703 507 6 vss
port 1 nsew
rlabel locali s 4134 474 4203 507 6 vss
port 1 nsew
rlabel locali s 3634 474 3703 507 6 vss
port 1 nsew
rlabel locali s 3134 474 3203 507 6 vss
port 1 nsew
rlabel locali s 2634 474 2703 507 6 vss
port 1 nsew
rlabel locali s 2134 474 2203 507 6 vss
port 1 nsew
rlabel locali s 1634 474 1703 507 6 vss
port 1 nsew
rlabel locali s 1134 474 1203 507 6 vss
port 1 nsew
rlabel locali s 634 474 703 507 6 vss
port 1 nsew
rlabel locali s 5044 606 5061 710 6 vss
port 1 nsew
rlabel locali s 4544 606 4561 710 6 vss
port 1 nsew
rlabel locali s 4044 606 4061 710 6 vss
port 1 nsew
rlabel locali s 3544 606 3561 710 6 vss
port 1 nsew
rlabel locali s 3044 606 3061 710 6 vss
port 1 nsew
rlabel locali s 2544 606 2561 710 6 vss
port 1 nsew
rlabel locali s 2044 606 2061 710 6 vss
port 1 nsew
rlabel locali s 1544 606 1561 710 6 vss
port 1 nsew
rlabel locali s 1044 606 1061 710 6 vss
port 1 nsew
rlabel locali s 544 606 561 710 6 vss
port 1 nsew
rlabel locali s 5044 856 5061 960 6 vss
port 1 nsew
rlabel locali s 4544 856 4561 960 6 vss
port 1 nsew
rlabel locali s 4044 856 4061 960 6 vss
port 1 nsew
rlabel locali s 3544 856 3561 960 6 vss
port 1 nsew
rlabel locali s 3044 856 3061 960 6 vss
port 1 nsew
rlabel locali s 2544 856 2561 960 6 vss
port 1 nsew
rlabel locali s 2044 856 2061 960 6 vss
port 1 nsew
rlabel locali s 1544 856 1561 960 6 vss
port 1 nsew
rlabel locali s 1044 856 1061 960 6 vss
port 1 nsew
rlabel locali s 544 856 561 960 6 vss
port 1 nsew
rlabel locali s 5135 1042 5204 1075 6 vss
port 1 nsew
rlabel locali s 4635 1042 4704 1075 6 vss
port 1 nsew
rlabel locali s 4135 1042 4204 1075 6 vss
port 1 nsew
rlabel locali s 3635 1042 3704 1075 6 vss
port 1 nsew
rlabel locali s 3135 1042 3204 1075 6 vss
port 1 nsew
rlabel locali s 2635 1042 2704 1075 6 vss
port 1 nsew
rlabel locali s 2135 1042 2204 1075 6 vss
port 1 nsew
rlabel locali s 1635 1042 1704 1075 6 vss
port 1 nsew
rlabel locali s 1135 1042 1204 1075 6 vss
port 1 nsew
rlabel locali s 635 1042 704 1075 6 vss
port 1 nsew
rlabel locali s 10541 3740 10574 3810 6 vss
port 1 nsew
rlabel metal2 s 634 763 5214 805 6 bias
port 2 nsew
rlabel via1 s 5174 771 5200 797 6 bias
port 2 nsew
rlabel via1 s 5142 771 5168 797 6 bias
port 2 nsew
rlabel via1 s 4674 771 4700 797 6 bias
port 2 nsew
rlabel via1 s 4642 771 4668 797 6 bias
port 2 nsew
rlabel via1 s 4174 771 4200 797 6 bias
port 2 nsew
rlabel via1 s 4142 771 4168 797 6 bias
port 2 nsew
rlabel via1 s 3674 771 3700 797 6 bias
port 2 nsew
rlabel via1 s 3642 771 3668 797 6 bias
port 2 nsew
rlabel via1 s 3174 771 3200 797 6 bias
port 2 nsew
rlabel via1 s 3142 771 3168 797 6 bias
port 2 nsew
rlabel via1 s 2674 771 2700 797 6 bias
port 2 nsew
rlabel via1 s 2642 771 2668 797 6 bias
port 2 nsew
rlabel via1 s 2174 771 2200 797 6 bias
port 2 nsew
rlabel via1 s 2142 771 2168 797 6 bias
port 2 nsew
rlabel via1 s 1674 771 1700 797 6 bias
port 2 nsew
rlabel via1 s 1642 771 1668 797 6 bias
port 2 nsew
rlabel via1 s 1174 771 1200 797 6 bias
port 2 nsew
rlabel via1 s 1142 771 1168 797 6 bias
port 2 nsew
rlabel via1 s 674 771 700 797 6 bias
port 2 nsew
rlabel via1 s 642 771 668 797 6 bias
port 2 nsew
rlabel metal1 s 5069 569 5265 592 6 bias
port 2 nsew
rlabel metal1 s 4569 569 4765 592 6 bias
port 2 nsew
rlabel metal1 s 4069 569 4265 592 6 bias
port 2 nsew
rlabel metal1 s 3569 569 3765 592 6 bias
port 2 nsew
rlabel metal1 s 3069 569 3265 592 6 bias
port 2 nsew
rlabel metal1 s 2569 569 2765 592 6 bias
port 2 nsew
rlabel metal1 s 2069 569 2265 592 6 bias
port 2 nsew
rlabel metal1 s 1569 569 1765 592 6 bias
port 2 nsew
rlabel metal1 s 1069 569 1265 592 6 bias
port 2 nsew
rlabel metal1 s 793 430 856 608 6 bias
port 2 nsew
rlabel metal1 s 569 569 765 592 6 bias
port 2 nsew
rlabel metal1 s 770 608 856 708 6 bias
port 2 nsew
rlabel metal1 s 5069 724 5265 842 6 bias
port 2 nsew
rlabel metal1 s 4569 724 4765 842 6 bias
port 2 nsew
rlabel metal1 s 4069 724 4265 842 6 bias
port 2 nsew
rlabel metal1 s 3569 724 3765 842 6 bias
port 2 nsew
rlabel metal1 s 3069 724 3265 842 6 bias
port 2 nsew
rlabel metal1 s 2569 724 2765 842 6 bias
port 2 nsew
rlabel metal1 s 2069 724 2265 842 6 bias
port 2 nsew
rlabel metal1 s 1569 724 1765 842 6 bias
port 2 nsew
rlabel metal1 s 1069 724 1265 842 6 bias
port 2 nsew
rlabel metal1 s 793 708 856 747 6 bias
port 2 nsew
rlabel metal1 s 569 724 765 747 6 bias
port 2 nsew
rlabel metal1 s 569 747 856 819 6 bias
port 2 nsew
rlabel metal1 s 793 819 856 858 6 bias
port 2 nsew
rlabel metal1 s 569 819 765 842 6 bias
port 2 nsew
rlabel metal1 s 770 858 856 958 6 bias
port 2 nsew
rlabel metal1 s 5069 974 5265 997 6 bias
port 2 nsew
rlabel metal1 s 4569 974 4765 997 6 bias
port 2 nsew
rlabel metal1 s 4069 974 4265 997 6 bias
port 2 nsew
rlabel metal1 s 3569 974 3765 997 6 bias
port 2 nsew
rlabel metal1 s 3069 974 3265 997 6 bias
port 2 nsew
rlabel metal1 s 2569 974 2765 997 6 bias
port 2 nsew
rlabel metal1 s 2069 974 2265 997 6 bias
port 2 nsew
rlabel metal1 s 1569 974 1765 997 6 bias
port 2 nsew
rlabel metal1 s 1069 974 1265 997 6 bias
port 2 nsew
rlabel metal1 s 793 958 856 1144 6 bias
port 2 nsew
rlabel metal1 s 569 974 765 997 6 bias
port 2 nsew
rlabel metal1 s -4600 1144 856 1206 4 bias
port 2 nsew
rlabel locali s 5067 572 5267 589 6 bias
port 2 nsew
rlabel locali s 4567 572 4767 589 6 bias
port 2 nsew
rlabel locali s 4067 572 4267 589 6 bias
port 2 nsew
rlabel locali s 3567 572 3767 589 6 bias
port 2 nsew
rlabel locali s 3067 572 3267 589 6 bias
port 2 nsew
rlabel locali s 2567 572 2767 589 6 bias
port 2 nsew
rlabel locali s 2067 572 2267 589 6 bias
port 2 nsew
rlabel locali s 1567 572 1767 589 6 bias
port 2 nsew
rlabel locali s 1067 572 1267 589 6 bias
port 2 nsew
rlabel locali s 567 572 767 589 6 bias
port 2 nsew
rlabel locali s 773 606 790 710 6 bias
port 2 nsew
rlabel locali s 5067 727 5267 744 6 bias
port 2 nsew
rlabel locali s 4567 727 4767 744 6 bias
port 2 nsew
rlabel locali s 4067 727 4267 744 6 bias
port 2 nsew
rlabel locali s 3567 727 3767 744 6 bias
port 2 nsew
rlabel locali s 3067 727 3267 744 6 bias
port 2 nsew
rlabel locali s 2567 727 2767 744 6 bias
port 2 nsew
rlabel locali s 2067 727 2267 744 6 bias
port 2 nsew
rlabel locali s 1567 727 1767 744 6 bias
port 2 nsew
rlabel locali s 1067 727 1267 744 6 bias
port 2 nsew
rlabel locali s 567 727 767 744 6 bias
port 2 nsew
rlabel locali s 5067 822 5267 839 6 bias
port 2 nsew
rlabel locali s 4567 822 4767 839 6 bias
port 2 nsew
rlabel locali s 4067 822 4267 839 6 bias
port 2 nsew
rlabel locali s 3567 822 3767 839 6 bias
port 2 nsew
rlabel locali s 3067 822 3267 839 6 bias
port 2 nsew
rlabel locali s 2567 822 2767 839 6 bias
port 2 nsew
rlabel locali s 2067 822 2267 839 6 bias
port 2 nsew
rlabel locali s 1567 822 1767 839 6 bias
port 2 nsew
rlabel locali s 1067 822 1267 839 6 bias
port 2 nsew
rlabel locali s 567 822 767 839 6 bias
port 2 nsew
rlabel locali s 773 856 790 960 6 bias
port 2 nsew
rlabel locali s 5067 977 5267 994 6 bias
port 2 nsew
rlabel locali s 4567 977 4767 994 6 bias
port 2 nsew
rlabel locali s 4067 977 4267 994 6 bias
port 2 nsew
rlabel locali s 3567 977 3767 994 6 bias
port 2 nsew
rlabel locali s 3067 977 3267 994 6 bias
port 2 nsew
rlabel locali s 2567 977 2767 994 6 bias
port 2 nsew
rlabel locali s 2067 977 2267 994 6 bias
port 2 nsew
rlabel locali s 1567 977 1767 994 6 bias
port 2 nsew
rlabel locali s 1067 977 1267 994 6 bias
port 2 nsew
rlabel locali s 567 977 767 994 6 bias
port 2 nsew
rlabel metal1 s 8929 2710 9159 2762 6 vdd
port 3 nsew
rlabel metal1 s 8479 2710 8709 2762 6 vdd
port 3 nsew
rlabel metal1 s 8029 2710 8259 2762 6 vdd
port 3 nsew
rlabel metal1 s 7579 2710 7809 2762 6 vdd
port 3 nsew
rlabel metal1 s 7129 2710 7359 2762 6 vdd
port 3 nsew
rlabel metal1 s 6679 2710 6909 2762 6 vdd
port 3 nsew
rlabel metal1 s 6229 2710 6459 2762 6 vdd
port 3 nsew
rlabel metal1 s 5779 2710 6009 2762 6 vdd
port 3 nsew
rlabel metal1 s 8929 2762 8995 2855 6 vdd
port 3 nsew
rlabel metal1 s 8479 2762 8545 2855 6 vdd
port 3 nsew
rlabel metal1 s 8029 2762 8095 2855 6 vdd
port 3 nsew
rlabel metal1 s 7579 2762 7645 2855 6 vdd
port 3 nsew
rlabel metal1 s 7129 2762 7195 2855 6 vdd
port 3 nsew
rlabel metal1 s 6679 2762 6745 2855 6 vdd
port 3 nsew
rlabel metal1 s 6229 2762 6295 2855 6 vdd
port 3 nsew
rlabel metal1 s 5779 2762 5845 2855 6 vdd
port 3 nsew
rlabel metal1 s 8929 2855 9018 3055 6 vdd
port 3 nsew
rlabel metal1 s 8479 2855 8568 3055 6 vdd
port 3 nsew
rlabel metal1 s 8029 2855 8118 3055 6 vdd
port 3 nsew
rlabel metal1 s 7579 2855 7668 3055 6 vdd
port 3 nsew
rlabel metal1 s 7129 2855 7218 3055 6 vdd
port 3 nsew
rlabel metal1 s 6679 2855 6768 3055 6 vdd
port 3 nsew
rlabel metal1 s 6229 2855 6318 3055 6 vdd
port 3 nsew
rlabel metal1 s 5779 2855 5868 3055 6 vdd
port 3 nsew
rlabel metal1 s 8929 3055 8995 3225 6 vdd
port 3 nsew
rlabel metal1 s 8479 3055 8545 3225 6 vdd
port 3 nsew
rlabel metal1 s 8029 3055 8095 3225 6 vdd
port 3 nsew
rlabel metal1 s 7579 3055 7645 3225 6 vdd
port 3 nsew
rlabel metal1 s 7129 3055 7195 3225 6 vdd
port 3 nsew
rlabel metal1 s 6679 3055 6745 3225 6 vdd
port 3 nsew
rlabel metal1 s 6229 3055 6295 3225 6 vdd
port 3 nsew
rlabel metal1 s 5779 3055 5845 3225 6 vdd
port 3 nsew
rlabel metal1 s 8929 3225 9018 3425 6 vdd
port 3 nsew
rlabel metal1 s 8479 3225 8568 3425 6 vdd
port 3 nsew
rlabel metal1 s 8029 3225 8118 3425 6 vdd
port 3 nsew
rlabel metal1 s 7579 3225 7668 3425 6 vdd
port 3 nsew
rlabel metal1 s 7129 3225 7218 3425 6 vdd
port 3 nsew
rlabel metal1 s 6679 3225 6768 3425 6 vdd
port 3 nsew
rlabel metal1 s 6229 3225 6318 3425 6 vdd
port 3 nsew
rlabel metal1 s 5779 3225 5868 3425 6 vdd
port 3 nsew
rlabel metal1 s 8929 3425 8995 3513 6 vdd
port 3 nsew
rlabel metal1 s 8479 3425 8545 3513 6 vdd
port 3 nsew
rlabel metal1 s 8029 3425 8095 3513 6 vdd
port 3 nsew
rlabel metal1 s 7579 3425 7645 3513 6 vdd
port 3 nsew
rlabel metal1 s 7129 3425 7195 3513 6 vdd
port 3 nsew
rlabel metal1 s 6679 3425 6745 3513 6 vdd
port 3 nsew
rlabel metal1 s 6229 3425 6295 3513 6 vdd
port 3 nsew
rlabel metal1 s 5779 3425 5845 3513 6 vdd
port 3 nsew
rlabel metal1 s 8929 3513 9159 3565 6 vdd
port 3 nsew
rlabel metal1 s 8479 3513 8709 3565 6 vdd
port 3 nsew
rlabel metal1 s 8029 3513 8259 3565 6 vdd
port 3 nsew
rlabel metal1 s 7579 3513 7809 3565 6 vdd
port 3 nsew
rlabel metal1 s 7129 3513 7359 3565 6 vdd
port 3 nsew
rlabel metal1 s 6679 3513 6909 3565 6 vdd
port 3 nsew
rlabel metal1 s 6229 3513 6459 3565 6 vdd
port 3 nsew
rlabel metal1 s 5779 3513 6009 3565 6 vdd
port 3 nsew
rlabel metal1 s 8929 3565 8995 3646 6 vdd
port 3 nsew
rlabel metal1 s 8479 3565 8545 3646 6 vdd
port 3 nsew
rlabel metal1 s 8029 3565 8095 3646 6 vdd
port 3 nsew
rlabel metal1 s 7579 3565 7645 3646 6 vdd
port 3 nsew
rlabel metal1 s 7129 3565 7195 3646 6 vdd
port 3 nsew
rlabel metal1 s 6679 3565 6745 3646 6 vdd
port 3 nsew
rlabel metal1 s 6229 3565 6295 3646 6 vdd
port 3 nsew
rlabel metal1 s 5779 3565 5845 3646 6 vdd
port 3 nsew
rlabel metal1 s 1420 3540 1650 3592 6 vdd
port 3 nsew
rlabel metal1 s 920 3540 1150 3592 6 vdd
port 3 nsew
rlabel metal1 s 2063 3646 8995 3737 6 vdd
port 3 nsew
rlabel metal1 s 1420 3592 1486 3685 6 vdd
port 3 nsew
rlabel metal1 s 920 3592 986 3685 6 vdd
port 3 nsew
rlabel metal1 s 2063 3737 2133 4476 6 vdd
port 3 nsew
rlabel metal1 s 1420 3685 1509 3885 6 vdd
port 3 nsew
rlabel metal1 s 920 3685 1009 3885 6 vdd
port 3 nsew
rlabel metal1 s 1420 3885 1486 4055 6 vdd
port 3 nsew
rlabel metal1 s 920 3885 986 4055 6 vdd
port 3 nsew
rlabel metal1 s 1420 4055 1509 4255 6 vdd
port 3 nsew
rlabel metal1 s 920 4055 1009 4255 6 vdd
port 3 nsew
rlabel metal1 s 1420 4255 1486 4343 6 vdd
port 3 nsew
rlabel metal1 s 920 4255 986 4343 6 vdd
port 3 nsew
rlabel metal1 s 1420 4343 1650 4395 6 vdd
port 3 nsew
rlabel metal1 s 920 4343 1150 4395 6 vdd
port 3 nsew
rlabel metal1 s 1420 4395 1486 4476 6 vdd
port 3 nsew
rlabel metal1 s 920 4395 986 4476 6 vdd
port 3 nsew
rlabel metal1 s -4600 4476 2133 4535 4 vdd
port 3 nsew
rlabel locali s 9083 2720 9152 2753 6 vdd
port 3 nsew
rlabel locali s 8633 2720 8702 2753 6 vdd
port 3 nsew
rlabel locali s 8183 2720 8252 2753 6 vdd
port 3 nsew
rlabel locali s 7733 2720 7802 2753 6 vdd
port 3 nsew
rlabel locali s 7283 2720 7352 2753 6 vdd
port 3 nsew
rlabel locali s 6833 2720 6902 2753 6 vdd
port 3 nsew
rlabel locali s 6383 2720 6452 2753 6 vdd
port 3 nsew
rlabel locali s 5933 2720 6002 2753 6 vdd
port 3 nsew
rlabel locali s 8998 2853 9015 3057 6 vdd
port 3 nsew
rlabel locali s 8548 2853 8565 3057 6 vdd
port 3 nsew
rlabel locali s 8098 2853 8115 3057 6 vdd
port 3 nsew
rlabel locali s 7648 2853 7665 3057 6 vdd
port 3 nsew
rlabel locali s 7198 2853 7215 3057 6 vdd
port 3 nsew
rlabel locali s 6748 2853 6765 3057 6 vdd
port 3 nsew
rlabel locali s 6298 2853 6315 3057 6 vdd
port 3 nsew
rlabel locali s 5848 2853 5865 3057 6 vdd
port 3 nsew
rlabel locali s 8998 3223 9015 3427 6 vdd
port 3 nsew
rlabel locali s 8548 3223 8565 3427 6 vdd
port 3 nsew
rlabel locali s 8098 3223 8115 3427 6 vdd
port 3 nsew
rlabel locali s 7648 3223 7665 3427 6 vdd
port 3 nsew
rlabel locali s 7198 3223 7215 3427 6 vdd
port 3 nsew
rlabel locali s 6748 3223 6765 3427 6 vdd
port 3 nsew
rlabel locali s 6298 3223 6315 3427 6 vdd
port 3 nsew
rlabel locali s 5848 3223 5865 3427 6 vdd
port 3 nsew
rlabel locali s 9085 3522 9154 3555 6 vdd
port 3 nsew
rlabel locali s 8635 3522 8704 3555 6 vdd
port 3 nsew
rlabel locali s 8185 3522 8254 3555 6 vdd
port 3 nsew
rlabel locali s 7735 3522 7804 3555 6 vdd
port 3 nsew
rlabel locali s 7285 3522 7354 3555 6 vdd
port 3 nsew
rlabel locali s 6835 3522 6904 3555 6 vdd
port 3 nsew
rlabel locali s 6385 3522 6454 3555 6 vdd
port 3 nsew
rlabel locali s 5935 3522 6004 3555 6 vdd
port 3 nsew
rlabel locali s 1574 3550 1643 3583 6 vdd
port 3 nsew
rlabel locali s 1074 3550 1143 3583 6 vdd
port 3 nsew
rlabel locali s 1489 3683 1506 3887 6 vdd
port 3 nsew
rlabel locali s 989 3683 1006 3887 6 vdd
port 3 nsew
rlabel locali s 1489 4053 1506 4257 6 vdd
port 3 nsew
rlabel locali s 989 4053 1006 4257 6 vdd
port 3 nsew
rlabel locali s 1576 4352 1645 4385 6 vdd
port 3 nsew
rlabel locali s 1076 4352 1145 4385 6 vdd
port 3 nsew
rlabel metal1 s 5293 430 5356 608 6 out
port 4 nsew
rlabel metal1 s 4793 430 4856 608 6 out
port 4 nsew
rlabel metal1 s 4293 430 4356 608 6 out
port 4 nsew
rlabel metal1 s 3793 430 3856 608 6 out
port 4 nsew
rlabel metal1 s 3293 430 3356 608 6 out
port 4 nsew
rlabel metal1 s 2793 430 2856 608 6 out
port 4 nsew
rlabel metal1 s 2293 430 2356 608 6 out
port 4 nsew
rlabel metal1 s 1793 430 1856 608 6 out
port 4 nsew
rlabel metal1 s 5270 608 5356 708 6 out
port 4 nsew
rlabel metal1 s 4770 608 4856 708 6 out
port 4 nsew
rlabel metal1 s 4270 608 4356 708 6 out
port 4 nsew
rlabel metal1 s 3770 608 3856 708 6 out
port 4 nsew
rlabel metal1 s 3270 608 3356 708 6 out
port 4 nsew
rlabel metal1 s 2770 608 2856 708 6 out
port 4 nsew
rlabel metal1 s 2270 608 2356 708 6 out
port 4 nsew
rlabel metal1 s 1770 608 1856 708 6 out
port 4 nsew
rlabel metal1 s 5293 708 5356 858 6 out
port 4 nsew
rlabel metal1 s 4793 708 4856 858 6 out
port 4 nsew
rlabel metal1 s 4293 708 4356 858 6 out
port 4 nsew
rlabel metal1 s 3793 708 3856 858 6 out
port 4 nsew
rlabel metal1 s 3293 708 3356 858 6 out
port 4 nsew
rlabel metal1 s 2793 708 2856 858 6 out
port 4 nsew
rlabel metal1 s 2293 708 2356 858 6 out
port 4 nsew
rlabel metal1 s 1793 708 1856 858 6 out
port 4 nsew
rlabel metal1 s 5270 858 5356 958 6 out
port 4 nsew
rlabel metal1 s 4770 858 4856 958 6 out
port 4 nsew
rlabel metal1 s 4270 858 4356 958 6 out
port 4 nsew
rlabel metal1 s 3770 858 3856 958 6 out
port 4 nsew
rlabel metal1 s 3270 858 3356 958 6 out
port 4 nsew
rlabel metal1 s 2770 858 2856 958 6 out
port 4 nsew
rlabel metal1 s 2270 858 2356 958 6 out
port 4 nsew
rlabel metal1 s 1770 858 1856 958 6 out
port 4 nsew
rlabel metal1 s 5293 958 5356 1199 6 out
port 4 nsew
rlabel metal1 s 4793 958 4856 1199 6 out
port 4 nsew
rlabel metal1 s 4293 958 4356 1199 6 out
port 4 nsew
rlabel metal1 s 3793 958 3856 1199 6 out
port 4 nsew
rlabel metal1 s 3293 958 3356 1199 6 out
port 4 nsew
rlabel metal1 s 2793 958 2856 1199 6 out
port 4 nsew
rlabel metal1 s 2293 958 2356 1199 6 out
port 4 nsew
rlabel metal1 s 1793 958 1856 1199 6 out
port 4 nsew
rlabel metal1 s 1793 1199 6231 1260 6 out
port 4 nsew
rlabel metal1 s 6146 1260 6231 1870 6 out
port 4 nsew
rlabel metal1 s 6146 1870 16925 1988 6 out
port 4 nsew
rlabel metal1 s 10725 1988 10784 3242 6 out
port 4 nsew
rlabel metal1 s 6146 1988 6231 2532 6 out
port 4 nsew
rlabel metal1 s 6097 2532 9314 2625 6 out
port 4 nsew
rlabel metal1 s 9247 2625 9314 2855 6 out
port 4 nsew
rlabel metal1 s 8797 2625 8864 2855 6 out
port 4 nsew
rlabel metal1 s 8347 2625 8414 2855 6 out
port 4 nsew
rlabel metal1 s 7897 2625 7964 2855 6 out
port 4 nsew
rlabel metal1 s 7447 2625 7514 2855 6 out
port 4 nsew
rlabel metal1 s 6997 2625 7064 2855 6 out
port 4 nsew
rlabel metal1 s 6547 2625 6614 2855 6 out
port 4 nsew
rlabel metal1 s 6097 2625 6164 2855 6 out
port 4 nsew
rlabel metal1 s 9224 2855 9314 3055 6 out
port 4 nsew
rlabel metal1 s 8774 2855 8864 3055 6 out
port 4 nsew
rlabel metal1 s 8324 2855 8414 3055 6 out
port 4 nsew
rlabel metal1 s 7874 2855 7964 3055 6 out
port 4 nsew
rlabel metal1 s 7424 2855 7514 3055 6 out
port 4 nsew
rlabel metal1 s 6974 2855 7064 3055 6 out
port 4 nsew
rlabel metal1 s 6524 2855 6614 3055 6 out
port 4 nsew
rlabel metal1 s 6074 2855 6164 3055 6 out
port 4 nsew
rlabel metal1 s 9247 3055 9314 3225 6 out
port 4 nsew
rlabel metal1 s 8797 3055 8864 3225 6 out
port 4 nsew
rlabel metal1 s 8347 3055 8414 3225 6 out
port 4 nsew
rlabel metal1 s 7897 3055 7964 3225 6 out
port 4 nsew
rlabel metal1 s 7447 3055 7514 3225 6 out
port 4 nsew
rlabel metal1 s 6997 3055 7064 3225 6 out
port 4 nsew
rlabel metal1 s 6547 3055 6614 3225 6 out
port 4 nsew
rlabel metal1 s 6097 3055 6164 3225 6 out
port 4 nsew
rlabel metal1 s 9224 3225 9314 3425 6 out
port 4 nsew
rlabel metal1 s 8774 3225 8864 3425 6 out
port 4 nsew
rlabel metal1 s 8324 3225 8414 3425 6 out
port 4 nsew
rlabel metal1 s 7874 3225 7964 3425 6 out
port 4 nsew
rlabel metal1 s 7424 3225 7514 3425 6 out
port 4 nsew
rlabel metal1 s 6974 3225 7064 3425 6 out
port 4 nsew
rlabel metal1 s 6524 3225 6614 3425 6 out
port 4 nsew
rlabel metal1 s 6074 3225 6164 3425 6 out
port 4 nsew
rlabel metal1 s 9247 3425 9314 3490 6 out
port 4 nsew
rlabel metal1 s 8797 3425 8864 3490 6 out
port 4 nsew
rlabel metal1 s 8347 3425 8414 3490 6 out
port 4 nsew
rlabel metal1 s 7897 3425 7964 3490 6 out
port 4 nsew
rlabel metal1 s 7447 3425 7514 3490 6 out
port 4 nsew
rlabel metal1 s 6997 3425 7064 3490 6 out
port 4 nsew
rlabel metal1 s 6547 3425 6614 3490 6 out
port 4 nsew
rlabel metal1 s 6097 3425 6164 3490 6 out
port 4 nsew
rlabel locali s 5273 606 5290 710 6 out
port 4 nsew
rlabel locali s 4773 606 4790 710 6 out
port 4 nsew
rlabel locali s 4273 606 4290 710 6 out
port 4 nsew
rlabel locali s 3773 606 3790 710 6 out
port 4 nsew
rlabel locali s 3273 606 3290 710 6 out
port 4 nsew
rlabel locali s 2773 606 2790 710 6 out
port 4 nsew
rlabel locali s 2273 606 2290 710 6 out
port 4 nsew
rlabel locali s 1773 606 1790 710 6 out
port 4 nsew
rlabel locali s 5273 856 5290 960 6 out
port 4 nsew
rlabel locali s 4773 856 4790 960 6 out
port 4 nsew
rlabel locali s 4273 856 4290 960 6 out
port 4 nsew
rlabel locali s 3773 856 3790 960 6 out
port 4 nsew
rlabel locali s 3273 856 3290 960 6 out
port 4 nsew
rlabel locali s 2773 856 2790 960 6 out
port 4 nsew
rlabel locali s 2273 856 2290 960 6 out
port 4 nsew
rlabel locali s 1773 856 1790 960 6 out
port 4 nsew
rlabel locali s 10720 3028 10789 3244 6 out
port 4 nsew
rlabel locali s 9227 2853 9244 3057 6 out
port 4 nsew
rlabel locali s 8777 2853 8794 3057 6 out
port 4 nsew
rlabel locali s 8327 2853 8344 3057 6 out
port 4 nsew
rlabel locali s 7877 2853 7894 3057 6 out
port 4 nsew
rlabel locali s 7427 2853 7444 3057 6 out
port 4 nsew
rlabel locali s 6977 2853 6994 3057 6 out
port 4 nsew
rlabel locali s 6527 2853 6544 3057 6 out
port 4 nsew
rlabel locali s 6077 2853 6094 3057 6 out
port 4 nsew
rlabel locali s 9227 3223 9244 3427 6 out
port 4 nsew
rlabel locali s 8777 3223 8794 3427 6 out
port 4 nsew
rlabel locali s 8327 3223 8344 3427 6 out
port 4 nsew
rlabel locali s 7877 3223 7894 3427 6 out
port 4 nsew
rlabel locali s 7427 3223 7444 3427 6 out
port 4 nsew
rlabel locali s 6977 3223 6994 3427 6 out
port 4 nsew
rlabel locali s 6527 3223 6544 3427 6 out
port 4 nsew
rlabel locali s 6077 3223 6094 3427 6 out
port 4 nsew
rlabel metal2 s -4600 1707 1137 1750 4 in_n
port 5 nsew
rlabel via1 s 1100 1716 1126 1742 6 in_n
port 5 nsew
rlabel via1 s 1068 1716 1094 1742 6 in_n
port 5 nsew
rlabel via1 s 750 1716 776 1742 6 in_n
port 5 nsew
rlabel via1 s 718 1716 744 1742 6 in_n
port 5 nsew
rlabel via1 s 400 1716 426 1742 6 in_n
port 5 nsew
rlabel via1 s 368 1716 394 1742 6 in_n
port 5 nsew
rlabel via1 s 50 1716 76 1742 6 in_n
port 5 nsew
rlabel via1 s 18 1716 44 1742 6 in_n
port 5 nsew
rlabel via1 s -301 1716 -275 1742 4 in_n
port 5 nsew
rlabel via1 s -333 1716 -307 1742 4 in_n
port 5 nsew
rlabel via1 s -651 1716 -625 1742 4 in_n
port 5 nsew
rlabel via1 s -683 1716 -657 1742 4 in_n
port 5 nsew
rlabel via1 s -1001 1716 -975 1742 4 in_n
port 5 nsew
rlabel via1 s -1033 1716 -1007 1742 4 in_n
port 5 nsew
rlabel via1 s -1351 1716 -1325 1742 4 in_n
port 5 nsew
rlabel via1 s -1383 1716 -1357 1742 4 in_n
port 5 nsew
rlabel via1 s -1701 1716 -1675 1742 4 in_n
port 5 nsew
rlabel via1 s -1733 1716 -1707 1742 4 in_n
port 5 nsew
rlabel via1 s -2051 1716 -2025 1742 4 in_n
port 5 nsew
rlabel via1 s -2083 1716 -2057 1742 4 in_n
port 5 nsew
rlabel metal1 s 1048 1679 1144 1799 6 in_n
port 5 nsew
rlabel metal1 s 698 1679 794 1799 6 in_n
port 5 nsew
rlabel metal1 s 348 1679 444 1799 6 in_n
port 5 nsew
rlabel metal1 s -2 1679 94 1799 6 in_n
port 5 nsew
rlabel metal1 s -352 1679 -256 1799 4 in_n
port 5 nsew
rlabel metal1 s -702 1679 -606 1799 4 in_n
port 5 nsew
rlabel metal1 s -1052 1679 -956 1799 4 in_n
port 5 nsew
rlabel metal1 s -1402 1679 -1306 1799 4 in_n
port 5 nsew
rlabel metal1 s -1752 1679 -1656 1799 4 in_n
port 5 nsew
rlabel metal1 s -2102 1679 -2006 1799 4 in_n
port 5 nsew
rlabel metal1 s 1048 2831 1144 2854 6 in_n
port 5 nsew
rlabel metal1 s 698 2831 794 2854 6 in_n
port 5 nsew
rlabel metal1 s 348 2831 444 2854 6 in_n
port 5 nsew
rlabel metal1 s -2 2831 94 2854 6 in_n
port 5 nsew
rlabel metal1 s -352 2831 -256 2854 4 in_n
port 5 nsew
rlabel metal1 s -702 2831 -606 2854 4 in_n
port 5 nsew
rlabel metal1 s -1052 2831 -956 2854 4 in_n
port 5 nsew
rlabel metal1 s -1402 2831 -1306 2854 4 in_n
port 5 nsew
rlabel metal1 s -1752 2831 -1656 2854 4 in_n
port 5 nsew
rlabel metal1 s -2102 2831 -2006 2854 4 in_n
port 5 nsew
rlabel locali s 1046 1779 1146 1796 6 in_n
port 5 nsew
rlabel locali s 696 1779 796 1796 6 in_n
port 5 nsew
rlabel locali s 346 1779 446 1796 6 in_n
port 5 nsew
rlabel locali s -4 1779 96 1796 6 in_n
port 5 nsew
rlabel locali s -354 1779 -254 1796 4 in_n
port 5 nsew
rlabel locali s -704 1779 -604 1796 4 in_n
port 5 nsew
rlabel locali s -1054 1779 -954 1796 4 in_n
port 5 nsew
rlabel locali s -1404 1779 -1304 1796 4 in_n
port 5 nsew
rlabel locali s -1754 1779 -1654 1796 4 in_n
port 5 nsew
rlabel locali s -2104 1779 -2004 1796 4 in_n
port 5 nsew
rlabel locali s 1046 2834 1146 2851 6 in_n
port 5 nsew
rlabel locali s 696 2834 796 2851 6 in_n
port 5 nsew
rlabel locali s 346 2834 446 2851 6 in_n
port 5 nsew
rlabel locali s -4 2834 96 2851 6 in_n
port 5 nsew
rlabel locali s -354 2834 -254 2851 4 in_n
port 5 nsew
rlabel locali s -704 2834 -604 2851 4 in_n
port 5 nsew
rlabel locali s -1054 2834 -954 2851 4 in_n
port 5 nsew
rlabel locali s -1404 2834 -1304 2851 4 in_n
port 5 nsew
rlabel locali s -1754 2834 -1654 2851 4 in_n
port 5 nsew
rlabel locali s -2104 2834 -2004 2851 4 in_n
port 5 nsew
rlabel metal2 s 1910 1707 16925 1750 6 in_p
port 6 nsew
rlabel via1 s 5100 1716 5126 1742 6 in_p
port 6 nsew
rlabel via1 s 5068 1716 5094 1742 6 in_p
port 6 nsew
rlabel via1 s 4750 1716 4776 1742 6 in_p
port 6 nsew
rlabel via1 s 4718 1716 4744 1742 6 in_p
port 6 nsew
rlabel via1 s 4400 1716 4426 1742 6 in_p
port 6 nsew
rlabel via1 s 4368 1716 4394 1742 6 in_p
port 6 nsew
rlabel via1 s 4050 1716 4076 1742 6 in_p
port 6 nsew
rlabel via1 s 4018 1716 4044 1742 6 in_p
port 6 nsew
rlabel via1 s 3700 1716 3726 1742 6 in_p
port 6 nsew
rlabel via1 s 3668 1716 3694 1742 6 in_p
port 6 nsew
rlabel via1 s 3350 1716 3376 1742 6 in_p
port 6 nsew
rlabel via1 s 3318 1716 3344 1742 6 in_p
port 6 nsew
rlabel via1 s 3000 1716 3026 1742 6 in_p
port 6 nsew
rlabel via1 s 2968 1716 2994 1742 6 in_p
port 6 nsew
rlabel via1 s 2650 1716 2676 1742 6 in_p
port 6 nsew
rlabel via1 s 2618 1716 2644 1742 6 in_p
port 6 nsew
rlabel via1 s 2300 1716 2326 1742 6 in_p
port 6 nsew
rlabel via1 s 2268 1716 2294 1742 6 in_p
port 6 nsew
rlabel via1 s 1950 1716 1976 1742 6 in_p
port 6 nsew
rlabel via1 s 1918 1716 1944 1742 6 in_p
port 6 nsew
rlabel metal1 s 5048 1679 5144 1799 6 in_p
port 6 nsew
rlabel metal1 s 4698 1679 4794 1799 6 in_p
port 6 nsew
rlabel metal1 s 4348 1679 4444 1799 6 in_p
port 6 nsew
rlabel metal1 s 3998 1679 4094 1799 6 in_p
port 6 nsew
rlabel metal1 s 3648 1679 3744 1799 6 in_p
port 6 nsew
rlabel metal1 s 3298 1679 3394 1799 6 in_p
port 6 nsew
rlabel metal1 s 2948 1679 3044 1799 6 in_p
port 6 nsew
rlabel metal1 s 2598 1679 2694 1799 6 in_p
port 6 nsew
rlabel metal1 s 2248 1679 2344 1799 6 in_p
port 6 nsew
rlabel metal1 s 1898 1679 1994 1799 6 in_p
port 6 nsew
rlabel metal1 s 5048 2831 5144 2854 6 in_p
port 6 nsew
rlabel metal1 s 4698 2831 4794 2854 6 in_p
port 6 nsew
rlabel metal1 s 4348 2831 4444 2854 6 in_p
port 6 nsew
rlabel metal1 s 3998 2831 4094 2854 6 in_p
port 6 nsew
rlabel metal1 s 3648 2831 3744 2854 6 in_p
port 6 nsew
rlabel metal1 s 3298 2831 3394 2854 6 in_p
port 6 nsew
rlabel metal1 s 2948 2831 3044 2854 6 in_p
port 6 nsew
rlabel metal1 s 2598 2831 2694 2854 6 in_p
port 6 nsew
rlabel metal1 s 2248 2831 2344 2854 6 in_p
port 6 nsew
rlabel metal1 s 1898 2831 1994 2854 6 in_p
port 6 nsew
rlabel locali s 5046 1779 5146 1796 6 in_p
port 6 nsew
rlabel locali s 4696 1779 4796 1796 6 in_p
port 6 nsew
rlabel locali s 4346 1779 4446 1796 6 in_p
port 6 nsew
rlabel locali s 3996 1779 4096 1796 6 in_p
port 6 nsew
rlabel locali s 3646 1779 3746 1796 6 in_p
port 6 nsew
rlabel locali s 3296 1779 3396 1796 6 in_p
port 6 nsew
rlabel locali s 2946 1779 3046 1796 6 in_p
port 6 nsew
rlabel locali s 2596 1779 2696 1796 6 in_p
port 6 nsew
rlabel locali s 2246 1779 2346 1796 6 in_p
port 6 nsew
rlabel locali s 1896 1779 1996 1796 6 in_p
port 6 nsew
rlabel locali s 5046 2834 5146 2851 6 in_p
port 6 nsew
rlabel locali s 4696 2834 4796 2851 6 in_p
port 6 nsew
rlabel locali s 4346 2834 4446 2851 6 in_p
port 6 nsew
rlabel locali s 3996 2834 4096 2851 6 in_p
port 6 nsew
rlabel locali s 3646 2834 3746 2851 6 in_p
port 6 nsew
rlabel locali s 3296 2834 3396 2851 6 in_p
port 6 nsew
rlabel locali s 2946 2834 3046 2851 6 in_p
port 6 nsew
rlabel locali s 2596 2834 2696 2851 6 in_p
port 6 nsew
rlabel locali s 2246 2834 2346 2851 6 in_p
port 6 nsew
rlabel locali s 1896 2834 1996 2851 6 in_p
port 6 nsew
rlabel metal1 -4600 4476 -4570 4535 1 vdd
port 3 n
rlabel metal1 -4600 248 -4570 357 1 vss
port 1 n
rlabel metal1 -4600 1144 -4570 1206 1 bias
port 2 n
rlabel metal2 -4600 1707 -4570 1750 1 in_n
port 5 n
rlabel metal2 16895 1707 16925 1750 1 in_p
port 6 n
rlabel metal1 16895 1870 16925 1988 1 out
port 4 n
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX -9200 496 33850 17224
string GDS_FILE layout.gds
string GDS_START 424954
string GDS_END 428916
string LEFview TRUE
<< end >>
