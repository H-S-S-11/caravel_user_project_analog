magic
tech sky130A
timestamp 1633199623
<< error_p >>
rect -88 192 -58 195
rect 10 192 40 195
rect -88 174 -82 192
rect 10 174 16 192
rect -88 171 -58 174
rect 10 171 40 174
rect -39 36 -9 39
rect 59 36 89 39
rect -39 18 -33 36
rect 59 18 65 36
rect -39 15 -9 18
rect 59 15 89 18
rect -39 -19 -9 -16
rect 59 -19 89 -16
rect -39 -37 -33 -19
rect 59 -37 65 -19
rect -39 -40 -9 -37
rect 59 -40 89 -37
rect -88 -175 -58 -172
rect 10 -175 40 -172
rect -88 -193 -82 -175
rect 10 -193 16 -175
rect -88 -196 -58 -193
rect 10 -196 40 -193
<< dnwell >>
rect -291 -371 291 371
<< nsonos >>
rect -82 55 -64 155
rect -33 55 -15 155
rect 16 55 34 155
rect 65 55 83 155
rect -82 -156 -64 -56
rect -33 -156 -15 -56
rect 16 -156 34 -56
rect 65 -156 83 -56
<< ndiff >>
rect -112 149 -82 155
rect -112 61 -106 149
rect -88 61 -82 149
rect -112 55 -82 61
rect -64 149 -33 155
rect -64 61 -58 149
rect -39 61 -33 149
rect -64 55 -33 61
rect -15 149 16 155
rect -15 61 -9 149
rect 10 61 16 149
rect -15 55 16 61
rect 34 149 65 155
rect 34 61 40 149
rect 59 61 65 149
rect 34 55 65 61
rect 83 149 113 155
rect 83 61 89 149
rect 107 61 113 149
rect 83 55 113 61
rect -112 -62 -82 -56
rect -112 -150 -106 -62
rect -88 -150 -82 -62
rect -112 -156 -82 -150
rect -64 -62 -33 -56
rect -64 -150 -58 -62
rect -39 -150 -33 -62
rect -64 -156 -33 -150
rect -15 -62 16 -56
rect -15 -150 -9 -62
rect 10 -150 16 -62
rect -15 -156 16 -150
rect 34 -62 65 -56
rect 34 -150 40 -62
rect 59 -150 65 -62
rect 34 -156 65 -150
rect 83 -62 113 -56
rect 83 -150 89 -62
rect 107 -150 113 -62
rect 83 -156 113 -150
<< ndiffc >>
rect -106 61 -88 149
rect -58 61 -39 149
rect -9 61 10 149
rect 40 61 59 149
rect 89 61 107 149
rect -106 -150 -88 -62
rect -58 -150 -39 -62
rect -9 -150 10 -62
rect 40 -150 59 -62
rect 89 -150 107 -62
<< poly >>
rect -90 192 -56 200
rect -90 174 -82 192
rect -64 174 -56 192
rect -90 166 -56 174
rect 8 192 42 200
rect 8 174 16 192
rect 34 174 42 192
rect -82 155 -64 166
rect -33 155 -15 168
rect 8 166 42 174
rect 16 155 34 166
rect 65 155 83 168
rect -82 42 -64 55
rect -33 44 -15 55
rect -41 36 -7 44
rect 16 42 34 55
rect 65 44 83 55
rect -41 18 -33 36
rect -15 18 -7 36
rect -41 10 -7 18
rect 57 36 91 44
rect 57 18 65 36
rect 83 18 91 36
rect 57 10 91 18
rect -41 -19 -7 -11
rect -41 -37 -33 -19
rect -15 -37 -7 -19
rect -82 -56 -64 -43
rect -41 -45 -7 -37
rect 57 -19 91 -11
rect 57 -37 65 -19
rect 83 -37 91 -19
rect -33 -56 -15 -45
rect 16 -56 34 -43
rect 57 -45 91 -37
rect 65 -56 83 -45
rect -82 -167 -64 -156
rect -90 -175 -56 -167
rect -33 -169 -15 -156
rect 16 -167 34 -156
rect -90 -193 -82 -175
rect -64 -193 -56 -175
rect -90 -201 -56 -193
rect 8 -175 42 -167
rect 65 -169 83 -156
rect 8 -193 16 -175
rect 34 -193 42 -175
rect 8 -201 42 -193
<< polycont >>
rect -82 174 -64 192
rect 16 174 34 192
rect -33 18 -15 36
rect 65 18 83 36
rect -33 -37 -15 -19
rect 65 -37 83 -19
rect -82 -193 -64 -175
rect 16 -193 34 -175
<< locali >>
rect -90 174 -82 192
rect -64 174 -56 192
rect 8 174 16 192
rect 34 174 42 192
rect -106 149 -88 157
rect -106 53 -88 61
rect -58 149 -39 157
rect -58 53 -39 61
rect -9 149 10 157
rect -9 53 10 61
rect 40 149 59 157
rect 40 53 59 61
rect 89 149 107 157
rect 89 53 107 61
rect -41 18 -33 36
rect -15 18 -7 36
rect 57 18 65 36
rect 83 18 91 36
rect -41 -37 -33 -19
rect -15 -37 -7 -19
rect 57 -37 65 -19
rect 83 -37 91 -19
rect -106 -62 -88 -54
rect -106 -158 -88 -150
rect -58 -62 -39 -54
rect -58 -158 -39 -150
rect -9 -62 10 -54
rect -9 -158 10 -150
rect 40 -62 59 -54
rect 40 -158 59 -150
rect 89 -62 107 -54
rect 89 -158 107 -150
rect -90 -193 -82 -175
rect -64 -193 -56 -175
rect 8 -193 16 -175
rect 34 -193 42 -175
<< viali >>
rect -82 174 -64 192
rect 16 174 34 192
rect -106 61 -88 149
rect -58 61 -39 149
rect -9 61 10 149
rect 40 61 59 149
rect 89 61 107 149
rect -33 18 -15 36
rect 65 18 83 36
rect -33 -37 -15 -19
rect 65 -37 83 -19
rect -106 -150 -88 -62
rect -58 -150 -39 -62
rect -9 -150 10 -62
rect 40 -150 59 -62
rect 89 -150 107 -62
rect -82 -193 -64 -175
rect 16 -193 34 -175
<< metal1 >>
rect -88 192 -58 195
rect -88 174 -82 192
rect -64 174 -58 192
rect -88 171 -58 174
rect 10 192 40 195
rect 10 174 16 192
rect 34 174 40 192
rect 10 171 40 174
rect -109 149 -85 155
rect -109 61 -106 149
rect -88 61 -85 149
rect -109 55 -85 61
rect -61 149 -36 155
rect -61 61 -58 149
rect -39 61 -36 149
rect -61 55 -36 61
rect -12 149 13 155
rect -12 61 -9 149
rect 10 61 13 149
rect -12 55 13 61
rect 37 149 62 155
rect 37 61 40 149
rect 59 61 62 149
rect 37 55 62 61
rect 86 149 110 155
rect 86 61 89 149
rect 107 61 110 149
rect 86 55 110 61
rect -39 36 -9 39
rect -39 18 -33 36
rect -15 18 -9 36
rect -39 15 -9 18
rect 59 36 89 39
rect 59 18 65 36
rect 83 18 89 36
rect 59 15 89 18
rect -39 -19 -9 -16
rect -39 -37 -33 -19
rect -15 -37 -9 -19
rect -39 -40 -9 -37
rect 59 -19 89 -16
rect 59 -37 65 -19
rect 83 -37 89 -19
rect 59 -40 89 -37
rect -109 -62 -85 -56
rect -109 -150 -106 -62
rect -88 -150 -85 -62
rect -109 -156 -85 -150
rect -61 -62 -36 -56
rect -61 -150 -58 -62
rect -39 -150 -36 -62
rect -61 -156 -36 -150
rect -12 -62 13 -56
rect -12 -150 -9 -62
rect 10 -150 13 -62
rect -12 -156 13 -150
rect 37 -62 62 -56
rect 37 -150 40 -62
rect 59 -150 62 -62
rect 37 -156 62 -150
rect 86 -62 110 -56
rect 86 -150 89 -62
rect 107 -150 110 -62
rect 86 -156 110 -150
rect -88 -175 -58 -172
rect -88 -193 -82 -175
rect -64 -193 -58 -175
rect -88 -196 -58 -193
rect 10 -175 40 -172
rect 10 -193 16 -175
rect 34 -193 40 -175
rect 10 -196 40 -193
<< properties >>
string gencell sky130_fd_bs_flash__special_sonosfet_star
string parameters w 1 l 0.18 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
