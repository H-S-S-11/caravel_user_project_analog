magic
tech sky130A
timestamp 1634337368
<< dnwell >>
rect -1700 0 -500 800
<< pwell >>
rect -1600 100 -500 700
<< psubdiff >>
rect -2100 1000 1400 1200
rect -2100 900 -1900 1000
rect 1200 900 1400 1000
rect -650 510 -530 530
rect -650 240 -630 510
rect -550 240 -530 510
rect -650 220 -530 240
rect -2100 -400 -1900 -300
rect 1200 -400 1400 -300
rect -2100 -600 -1800 -400
rect 1100 -600 1400 -400
<< psubdiffcont >>
rect -2100 -300 -1900 900
rect -630 240 -550 510
rect 1200 -300 1400 900
rect -1800 -600 1100 -400
<< locali >>
rect -2150 900 -1850 950
rect -2150 -300 -2100 900
rect -1900 -300 -1850 900
rect -1470 390 -1380 1300
rect -1340 450 -1250 1300
rect -1210 390 -1120 1300
rect -1470 290 -1350 390
rect -1240 290 -1120 390
rect -1070 390 -980 1300
rect -940 450 -850 1300
rect -810 390 -720 1300
rect -440 800 -260 1300
rect -170 800 -50 1300
rect -20 800 40 1300
rect 70 800 110 1300
rect 150 800 190 1300
rect 240 850 280 1300
rect 310 850 350 1300
rect 240 800 285 850
rect 305 800 350 850
rect 390 800 430 1300
rect 470 800 510 1300
rect -1070 290 -950 390
rect -840 290 -720 390
rect -650 510 -530 530
rect -650 240 -630 510
rect -550 240 -530 510
rect 700 430 800 1300
rect 850 320 950 1300
rect -650 220 -530 240
rect -1400 160 -530 220
rect -650 -60 -530 160
rect -170 -60 -50 270
rect 700 220 950 320
rect 1150 900 1450 950
rect -650 -180 -50 -60
rect -2150 -350 -1850 -300
rect 1150 -300 1200 900
rect 1400 700 1450 900
rect 1400 -100 1600 700
rect 1400 -300 1450 -100
rect 1150 -350 1450 -300
rect -2150 -400 1450 -350
rect -2150 -600 -1800 -400
rect 1100 -600 1450 -400
rect -2150 -650 1450 -600
<< viali >>
rect 1600 -100 2400 700
<< metal1 >>
rect 1500 700 2700 800
rect 1500 -100 1600 700
rect 2400 -100 2700 700
rect 1500 -200 2700 -100
use sky130_fd_bs_flash__special_sonosfet_star_VH7TJW  sky130_fd_bs_flash__special_sonosfet_star_VH7TJW_0
timestamp 1633983039
transform 1 0 291 0 1 371
box -791 -371 409 429
use sky130_fd_bs_flash__special_sonosfet_star_JJF9VQ  sky130_fd_bs_flash__special_sonosfet_star_JJF9VQ_0
timestamp 1633982189
transform 1 0 -898 0 1 340
box -102 -140 108 150
use sky130_fd_bs_flash__special_sonosfet_star_JJF9VQ  sky130_fd_bs_flash__special_sonosfet_star_JJF9VQ_1
timestamp 1633982189
transform 1 0 -1298 0 1 340
box -102 -140 108 150
<< labels >>
rlabel metal1 2500 -200 2700 800 1 VGND
port 10 n
rlabel locali 70 1280 110 1300 1 SEL_BOT
port 11 n
rlabel locali 150 1280 190 1300 1 RA3
port 12 n
rlabel locali 240 1280 280 1300 1 RA2
port 13 n
rlabel locali 310 1280 350 1300 1 RA1
port 14 n
rlabel locali 390 1280 430 1300 1 RA0
port 15 n
rlabel locali 470 1280 510 1300 1 SEL_TOP
port 16 n
rlabel locali -20 1280 40 1300 1 FLASH_SOURCE
port 17 n
rlabel locali 700 1280 800 1300 1 BL0
port 18 n
rlabel locali 850 1280 950 1300 1 BL1
port 19 n
rlabel locali -170 1280 -50 1300 1 PWELL
port 2 n
rlabel locali -440 1280 -260 1300 1 DNWELL
port 1 n
rlabel locali -1470 1280 -1380 1300 1 FS0
port 6 n
rlabel locali -1340 1280 -1250 1300 1 FG0
port 4 n
rlabel locali -1210 1280 -1120 1300 1 FD0
port 7 n
rlabel locali -1070 1280 -980 1300 1 FS1
port 8 n
rlabel locali -940 1280 -850 1300 1 FG1
port 5 n
rlabel locali -810 1280 -720 1300 1 FD1
port 9 n
<< end >>
