magic
tech sky130A
magscale 1 2
timestamp 1636387338
<< nwell >>
rect 1886 6993 3562 8843
rect 11604 5333 18580 7183
<< pwell >>
rect 21047 7447 21181 7653
rect -4202 5841 -3996 5975
rect -3502 5841 -3296 5975
rect -2802 5841 -2596 5975
rect -2102 5841 -1896 5975
rect -1402 5841 -1196 5975
rect -702 5841 -496 5975
rect -2 5841 204 5975
rect 698 5841 904 5975
rect 1398 5841 1604 5975
rect 2098 5841 2304 5975
rect 3798 5841 4004 5975
rect 4498 5841 4704 5975
rect 5198 5841 5404 5975
rect 5898 5841 6104 5975
rect 6598 5841 6804 5975
rect 7298 5841 7504 5975
rect 7998 5841 8204 5975
rect 8698 5841 8904 5975
rect 9398 5841 9604 5975
rect 10098 5841 10304 5975
rect -4292 3604 -3924 5656
rect -3592 3604 -3224 5656
rect -2892 3604 -2524 5656
rect -2192 3604 -1824 5656
rect -1492 3604 -1124 5656
rect -792 3604 -424 5656
rect -92 3604 276 5656
rect 608 3604 976 5656
rect 1308 3604 1676 5656
rect 2008 3604 2376 5656
rect 3708 3604 4076 5656
rect 4408 3604 4776 5656
rect 5108 3604 5476 5656
rect 5808 3604 6176 5656
rect 6508 3604 6876 5656
rect 7208 3604 7576 5656
rect 7908 3604 8276 5656
rect 8608 3604 8976 5656
rect 9308 3604 9676 5656
rect 10008 3604 10376 5656
rect 1235 1942 1441 2184
rect 2235 1942 2441 2184
rect 3235 1942 3441 2184
rect 4235 1942 4441 2184
rect 5235 1942 5441 2184
rect 6235 1942 6441 2184
rect 7235 1942 7441 2184
rect 8235 1942 8441 2184
rect 9235 1942 9441 2184
rect 10235 1942 10441 2184
rect 1050 1690 1618 1942
rect 2050 1690 2618 1942
rect 3050 1690 3618 1942
rect 4050 1690 4618 1942
rect 5050 1690 5618 1942
rect 6050 1690 6618 1942
rect 7050 1690 7618 1942
rect 8050 1690 8618 1942
rect 9050 1690 9618 1942
rect 10050 1690 10618 1942
rect 1050 1190 1618 1442
rect 2050 1190 2618 1442
rect 3050 1190 3618 1442
rect 4050 1190 4618 1442
rect 5050 1190 5618 1442
rect 6050 1190 6618 1442
rect 7050 1190 7618 1442
rect 8050 1190 8618 1442
rect 9050 1190 9618 1442
rect 10050 1190 10618 1442
rect 1234 913 1440 1190
rect 2234 913 2440 1190
rect 3234 913 3440 1190
rect 4234 913 4440 1190
rect 5234 913 5440 1190
rect 6234 913 6440 1190
rect 7234 913 7440 1190
rect 8234 913 8440 1190
rect 9234 913 9440 1190
rect 10234 913 10440 1190
<< mvnmos >>
rect -4208 3630 -4008 5630
rect -3508 3630 -3308 5630
rect -2808 3630 -2608 5630
rect -2108 3630 -1908 5630
rect -1408 3630 -1208 5630
rect -708 3630 -508 5630
rect -8 3630 192 5630
rect 692 3630 892 5630
rect 1392 3630 1592 5630
rect 2092 3630 2292 5630
rect 3792 3630 3992 5630
rect 4492 3630 4692 5630
rect 5192 3630 5392 5630
rect 5892 3630 6092 5630
rect 6592 3630 6792 5630
rect 7292 3630 7492 5630
rect 7992 3630 8192 5630
rect 8692 3630 8892 5630
rect 9392 3630 9592 5630
rect 10092 3630 10292 5630
rect 1134 1716 1534 1916
rect 2134 1716 2534 1916
rect 3134 1716 3534 1916
rect 4134 1716 4534 1916
rect 5134 1716 5534 1916
rect 6134 1716 6534 1916
rect 7134 1716 7534 1916
rect 8134 1716 8534 1916
rect 9134 1716 9534 1916
rect 10134 1716 10534 1916
rect 1134 1216 1534 1416
rect 2134 1216 2534 1416
rect 3134 1216 3534 1416
rect 4134 1216 4534 1416
rect 5134 1216 5534 1416
rect 6134 1216 6534 1416
rect 7134 1216 7534 1416
rect 8134 1216 8534 1416
rect 9134 1216 9534 1416
rect 10134 1216 10534 1416
<< mvpmos >>
rect 2024 8109 2424 8509
rect 3024 8109 3424 8509
rect 2024 7369 2424 7769
rect 3024 7369 3424 7769
rect 11742 6449 12142 6849
rect 12642 6449 13042 6849
rect 13542 6449 13942 6849
rect 14442 6449 14842 6849
rect 15342 6449 15742 6849
rect 16242 6449 16642 6849
rect 17142 6449 17542 6849
rect 18042 6449 18442 6849
rect 11742 5709 12142 6109
rect 12642 5709 13042 6109
rect 13542 5709 13942 6109
rect 14442 5709 14842 6109
rect 15342 5709 15742 6109
rect 16242 5709 16642 6109
rect 17142 5709 17542 6109
rect 18042 5709 18442 6109
<< mvndiff >>
rect -4266 5599 -4208 5630
rect -4266 5565 -4254 5599
rect -4220 5565 -4208 5599
rect -4266 5531 -4208 5565
rect -4266 5497 -4254 5531
rect -4220 5497 -4208 5531
rect -4266 5463 -4208 5497
rect -4266 5429 -4254 5463
rect -4220 5429 -4208 5463
rect -4266 5395 -4208 5429
rect -4266 5361 -4254 5395
rect -4220 5361 -4208 5395
rect -4266 5327 -4208 5361
rect -4266 5293 -4254 5327
rect -4220 5293 -4208 5327
rect -4266 5259 -4208 5293
rect -4266 5225 -4254 5259
rect -4220 5225 -4208 5259
rect -4266 5191 -4208 5225
rect -4266 5157 -4254 5191
rect -4220 5157 -4208 5191
rect -4266 5123 -4208 5157
rect -4266 5089 -4254 5123
rect -4220 5089 -4208 5123
rect -4266 5055 -4208 5089
rect -4266 5021 -4254 5055
rect -4220 5021 -4208 5055
rect -4266 4987 -4208 5021
rect -4266 4953 -4254 4987
rect -4220 4953 -4208 4987
rect -4266 4919 -4208 4953
rect -4266 4885 -4254 4919
rect -4220 4885 -4208 4919
rect -4266 4851 -4208 4885
rect -4266 4817 -4254 4851
rect -4220 4817 -4208 4851
rect -4266 4783 -4208 4817
rect -4266 4749 -4254 4783
rect -4220 4749 -4208 4783
rect -4266 4715 -4208 4749
rect -4266 4681 -4254 4715
rect -4220 4681 -4208 4715
rect -4266 4647 -4208 4681
rect -4266 4613 -4254 4647
rect -4220 4613 -4208 4647
rect -4266 4579 -4208 4613
rect -4266 4545 -4254 4579
rect -4220 4545 -4208 4579
rect -4266 4511 -4208 4545
rect -4266 4477 -4254 4511
rect -4220 4477 -4208 4511
rect -4266 4443 -4208 4477
rect -4266 4409 -4254 4443
rect -4220 4409 -4208 4443
rect -4266 4375 -4208 4409
rect -4266 4341 -4254 4375
rect -4220 4341 -4208 4375
rect -4266 4307 -4208 4341
rect -4266 4273 -4254 4307
rect -4220 4273 -4208 4307
rect -4266 4239 -4208 4273
rect -4266 4205 -4254 4239
rect -4220 4205 -4208 4239
rect -4266 4171 -4208 4205
rect -4266 4137 -4254 4171
rect -4220 4137 -4208 4171
rect -4266 4103 -4208 4137
rect -4266 4069 -4254 4103
rect -4220 4069 -4208 4103
rect -4266 4035 -4208 4069
rect -4266 4001 -4254 4035
rect -4220 4001 -4208 4035
rect -4266 3967 -4208 4001
rect -4266 3933 -4254 3967
rect -4220 3933 -4208 3967
rect -4266 3899 -4208 3933
rect -4266 3865 -4254 3899
rect -4220 3865 -4208 3899
rect -4266 3831 -4208 3865
rect -4266 3797 -4254 3831
rect -4220 3797 -4208 3831
rect -4266 3763 -4208 3797
rect -4266 3729 -4254 3763
rect -4220 3729 -4208 3763
rect -4266 3695 -4208 3729
rect -4266 3661 -4254 3695
rect -4220 3661 -4208 3695
rect -4266 3630 -4208 3661
rect -4008 5599 -3950 5630
rect -4008 5565 -3996 5599
rect -3962 5565 -3950 5599
rect -4008 5531 -3950 5565
rect -4008 5497 -3996 5531
rect -3962 5497 -3950 5531
rect -4008 5463 -3950 5497
rect -4008 5429 -3996 5463
rect -3962 5429 -3950 5463
rect -4008 5395 -3950 5429
rect -4008 5361 -3996 5395
rect -3962 5361 -3950 5395
rect -4008 5327 -3950 5361
rect -4008 5293 -3996 5327
rect -3962 5293 -3950 5327
rect -4008 5259 -3950 5293
rect -4008 5225 -3996 5259
rect -3962 5225 -3950 5259
rect -4008 5191 -3950 5225
rect -4008 5157 -3996 5191
rect -3962 5157 -3950 5191
rect -4008 5123 -3950 5157
rect -4008 5089 -3996 5123
rect -3962 5089 -3950 5123
rect -4008 5055 -3950 5089
rect -4008 5021 -3996 5055
rect -3962 5021 -3950 5055
rect -4008 4987 -3950 5021
rect -4008 4953 -3996 4987
rect -3962 4953 -3950 4987
rect -4008 4919 -3950 4953
rect -4008 4885 -3996 4919
rect -3962 4885 -3950 4919
rect -4008 4851 -3950 4885
rect -4008 4817 -3996 4851
rect -3962 4817 -3950 4851
rect -4008 4783 -3950 4817
rect -4008 4749 -3996 4783
rect -3962 4749 -3950 4783
rect -4008 4715 -3950 4749
rect -4008 4681 -3996 4715
rect -3962 4681 -3950 4715
rect -4008 4647 -3950 4681
rect -4008 4613 -3996 4647
rect -3962 4613 -3950 4647
rect -4008 4579 -3950 4613
rect -4008 4545 -3996 4579
rect -3962 4545 -3950 4579
rect -4008 4511 -3950 4545
rect -4008 4477 -3996 4511
rect -3962 4477 -3950 4511
rect -4008 4443 -3950 4477
rect -4008 4409 -3996 4443
rect -3962 4409 -3950 4443
rect -4008 4375 -3950 4409
rect -4008 4341 -3996 4375
rect -3962 4341 -3950 4375
rect -4008 4307 -3950 4341
rect -4008 4273 -3996 4307
rect -3962 4273 -3950 4307
rect -4008 4239 -3950 4273
rect -4008 4205 -3996 4239
rect -3962 4205 -3950 4239
rect -4008 4171 -3950 4205
rect -4008 4137 -3996 4171
rect -3962 4137 -3950 4171
rect -4008 4103 -3950 4137
rect -4008 4069 -3996 4103
rect -3962 4069 -3950 4103
rect -4008 4035 -3950 4069
rect -4008 4001 -3996 4035
rect -3962 4001 -3950 4035
rect -4008 3967 -3950 4001
rect -4008 3933 -3996 3967
rect -3962 3933 -3950 3967
rect -4008 3899 -3950 3933
rect -4008 3865 -3996 3899
rect -3962 3865 -3950 3899
rect -4008 3831 -3950 3865
rect -4008 3797 -3996 3831
rect -3962 3797 -3950 3831
rect -4008 3763 -3950 3797
rect -4008 3729 -3996 3763
rect -3962 3729 -3950 3763
rect -4008 3695 -3950 3729
rect -4008 3661 -3996 3695
rect -3962 3661 -3950 3695
rect -4008 3630 -3950 3661
rect -3566 5599 -3508 5630
rect -3566 5565 -3554 5599
rect -3520 5565 -3508 5599
rect -3566 5531 -3508 5565
rect -3566 5497 -3554 5531
rect -3520 5497 -3508 5531
rect -3566 5463 -3508 5497
rect -3566 5429 -3554 5463
rect -3520 5429 -3508 5463
rect -3566 5395 -3508 5429
rect -3566 5361 -3554 5395
rect -3520 5361 -3508 5395
rect -3566 5327 -3508 5361
rect -3566 5293 -3554 5327
rect -3520 5293 -3508 5327
rect -3566 5259 -3508 5293
rect -3566 5225 -3554 5259
rect -3520 5225 -3508 5259
rect -3566 5191 -3508 5225
rect -3566 5157 -3554 5191
rect -3520 5157 -3508 5191
rect -3566 5123 -3508 5157
rect -3566 5089 -3554 5123
rect -3520 5089 -3508 5123
rect -3566 5055 -3508 5089
rect -3566 5021 -3554 5055
rect -3520 5021 -3508 5055
rect -3566 4987 -3508 5021
rect -3566 4953 -3554 4987
rect -3520 4953 -3508 4987
rect -3566 4919 -3508 4953
rect -3566 4885 -3554 4919
rect -3520 4885 -3508 4919
rect -3566 4851 -3508 4885
rect -3566 4817 -3554 4851
rect -3520 4817 -3508 4851
rect -3566 4783 -3508 4817
rect -3566 4749 -3554 4783
rect -3520 4749 -3508 4783
rect -3566 4715 -3508 4749
rect -3566 4681 -3554 4715
rect -3520 4681 -3508 4715
rect -3566 4647 -3508 4681
rect -3566 4613 -3554 4647
rect -3520 4613 -3508 4647
rect -3566 4579 -3508 4613
rect -3566 4545 -3554 4579
rect -3520 4545 -3508 4579
rect -3566 4511 -3508 4545
rect -3566 4477 -3554 4511
rect -3520 4477 -3508 4511
rect -3566 4443 -3508 4477
rect -3566 4409 -3554 4443
rect -3520 4409 -3508 4443
rect -3566 4375 -3508 4409
rect -3566 4341 -3554 4375
rect -3520 4341 -3508 4375
rect -3566 4307 -3508 4341
rect -3566 4273 -3554 4307
rect -3520 4273 -3508 4307
rect -3566 4239 -3508 4273
rect -3566 4205 -3554 4239
rect -3520 4205 -3508 4239
rect -3566 4171 -3508 4205
rect -3566 4137 -3554 4171
rect -3520 4137 -3508 4171
rect -3566 4103 -3508 4137
rect -3566 4069 -3554 4103
rect -3520 4069 -3508 4103
rect -3566 4035 -3508 4069
rect -3566 4001 -3554 4035
rect -3520 4001 -3508 4035
rect -3566 3967 -3508 4001
rect -3566 3933 -3554 3967
rect -3520 3933 -3508 3967
rect -3566 3899 -3508 3933
rect -3566 3865 -3554 3899
rect -3520 3865 -3508 3899
rect -3566 3831 -3508 3865
rect -3566 3797 -3554 3831
rect -3520 3797 -3508 3831
rect -3566 3763 -3508 3797
rect -3566 3729 -3554 3763
rect -3520 3729 -3508 3763
rect -3566 3695 -3508 3729
rect -3566 3661 -3554 3695
rect -3520 3661 -3508 3695
rect -3566 3630 -3508 3661
rect -3308 5599 -3250 5630
rect -3308 5565 -3296 5599
rect -3262 5565 -3250 5599
rect -3308 5531 -3250 5565
rect -3308 5497 -3296 5531
rect -3262 5497 -3250 5531
rect -3308 5463 -3250 5497
rect -3308 5429 -3296 5463
rect -3262 5429 -3250 5463
rect -3308 5395 -3250 5429
rect -3308 5361 -3296 5395
rect -3262 5361 -3250 5395
rect -3308 5327 -3250 5361
rect -3308 5293 -3296 5327
rect -3262 5293 -3250 5327
rect -3308 5259 -3250 5293
rect -3308 5225 -3296 5259
rect -3262 5225 -3250 5259
rect -3308 5191 -3250 5225
rect -3308 5157 -3296 5191
rect -3262 5157 -3250 5191
rect -3308 5123 -3250 5157
rect -3308 5089 -3296 5123
rect -3262 5089 -3250 5123
rect -3308 5055 -3250 5089
rect -3308 5021 -3296 5055
rect -3262 5021 -3250 5055
rect -3308 4987 -3250 5021
rect -3308 4953 -3296 4987
rect -3262 4953 -3250 4987
rect -3308 4919 -3250 4953
rect -3308 4885 -3296 4919
rect -3262 4885 -3250 4919
rect -3308 4851 -3250 4885
rect -3308 4817 -3296 4851
rect -3262 4817 -3250 4851
rect -3308 4783 -3250 4817
rect -3308 4749 -3296 4783
rect -3262 4749 -3250 4783
rect -3308 4715 -3250 4749
rect -3308 4681 -3296 4715
rect -3262 4681 -3250 4715
rect -3308 4647 -3250 4681
rect -3308 4613 -3296 4647
rect -3262 4613 -3250 4647
rect -3308 4579 -3250 4613
rect -3308 4545 -3296 4579
rect -3262 4545 -3250 4579
rect -3308 4511 -3250 4545
rect -3308 4477 -3296 4511
rect -3262 4477 -3250 4511
rect -3308 4443 -3250 4477
rect -3308 4409 -3296 4443
rect -3262 4409 -3250 4443
rect -3308 4375 -3250 4409
rect -3308 4341 -3296 4375
rect -3262 4341 -3250 4375
rect -3308 4307 -3250 4341
rect -3308 4273 -3296 4307
rect -3262 4273 -3250 4307
rect -3308 4239 -3250 4273
rect -3308 4205 -3296 4239
rect -3262 4205 -3250 4239
rect -3308 4171 -3250 4205
rect -3308 4137 -3296 4171
rect -3262 4137 -3250 4171
rect -3308 4103 -3250 4137
rect -3308 4069 -3296 4103
rect -3262 4069 -3250 4103
rect -3308 4035 -3250 4069
rect -3308 4001 -3296 4035
rect -3262 4001 -3250 4035
rect -3308 3967 -3250 4001
rect -3308 3933 -3296 3967
rect -3262 3933 -3250 3967
rect -3308 3899 -3250 3933
rect -3308 3865 -3296 3899
rect -3262 3865 -3250 3899
rect -3308 3831 -3250 3865
rect -3308 3797 -3296 3831
rect -3262 3797 -3250 3831
rect -3308 3763 -3250 3797
rect -3308 3729 -3296 3763
rect -3262 3729 -3250 3763
rect -3308 3695 -3250 3729
rect -3308 3661 -3296 3695
rect -3262 3661 -3250 3695
rect -3308 3630 -3250 3661
rect -2866 5599 -2808 5630
rect -2866 5565 -2854 5599
rect -2820 5565 -2808 5599
rect -2866 5531 -2808 5565
rect -2866 5497 -2854 5531
rect -2820 5497 -2808 5531
rect -2866 5463 -2808 5497
rect -2866 5429 -2854 5463
rect -2820 5429 -2808 5463
rect -2866 5395 -2808 5429
rect -2866 5361 -2854 5395
rect -2820 5361 -2808 5395
rect -2866 5327 -2808 5361
rect -2866 5293 -2854 5327
rect -2820 5293 -2808 5327
rect -2866 5259 -2808 5293
rect -2866 5225 -2854 5259
rect -2820 5225 -2808 5259
rect -2866 5191 -2808 5225
rect -2866 5157 -2854 5191
rect -2820 5157 -2808 5191
rect -2866 5123 -2808 5157
rect -2866 5089 -2854 5123
rect -2820 5089 -2808 5123
rect -2866 5055 -2808 5089
rect -2866 5021 -2854 5055
rect -2820 5021 -2808 5055
rect -2866 4987 -2808 5021
rect -2866 4953 -2854 4987
rect -2820 4953 -2808 4987
rect -2866 4919 -2808 4953
rect -2866 4885 -2854 4919
rect -2820 4885 -2808 4919
rect -2866 4851 -2808 4885
rect -2866 4817 -2854 4851
rect -2820 4817 -2808 4851
rect -2866 4783 -2808 4817
rect -2866 4749 -2854 4783
rect -2820 4749 -2808 4783
rect -2866 4715 -2808 4749
rect -2866 4681 -2854 4715
rect -2820 4681 -2808 4715
rect -2866 4647 -2808 4681
rect -2866 4613 -2854 4647
rect -2820 4613 -2808 4647
rect -2866 4579 -2808 4613
rect -2866 4545 -2854 4579
rect -2820 4545 -2808 4579
rect -2866 4511 -2808 4545
rect -2866 4477 -2854 4511
rect -2820 4477 -2808 4511
rect -2866 4443 -2808 4477
rect -2866 4409 -2854 4443
rect -2820 4409 -2808 4443
rect -2866 4375 -2808 4409
rect -2866 4341 -2854 4375
rect -2820 4341 -2808 4375
rect -2866 4307 -2808 4341
rect -2866 4273 -2854 4307
rect -2820 4273 -2808 4307
rect -2866 4239 -2808 4273
rect -2866 4205 -2854 4239
rect -2820 4205 -2808 4239
rect -2866 4171 -2808 4205
rect -2866 4137 -2854 4171
rect -2820 4137 -2808 4171
rect -2866 4103 -2808 4137
rect -2866 4069 -2854 4103
rect -2820 4069 -2808 4103
rect -2866 4035 -2808 4069
rect -2866 4001 -2854 4035
rect -2820 4001 -2808 4035
rect -2866 3967 -2808 4001
rect -2866 3933 -2854 3967
rect -2820 3933 -2808 3967
rect -2866 3899 -2808 3933
rect -2866 3865 -2854 3899
rect -2820 3865 -2808 3899
rect -2866 3831 -2808 3865
rect -2866 3797 -2854 3831
rect -2820 3797 -2808 3831
rect -2866 3763 -2808 3797
rect -2866 3729 -2854 3763
rect -2820 3729 -2808 3763
rect -2866 3695 -2808 3729
rect -2866 3661 -2854 3695
rect -2820 3661 -2808 3695
rect -2866 3630 -2808 3661
rect -2608 5599 -2550 5630
rect -2608 5565 -2596 5599
rect -2562 5565 -2550 5599
rect -2608 5531 -2550 5565
rect -2608 5497 -2596 5531
rect -2562 5497 -2550 5531
rect -2608 5463 -2550 5497
rect -2608 5429 -2596 5463
rect -2562 5429 -2550 5463
rect -2608 5395 -2550 5429
rect -2608 5361 -2596 5395
rect -2562 5361 -2550 5395
rect -2608 5327 -2550 5361
rect -2608 5293 -2596 5327
rect -2562 5293 -2550 5327
rect -2608 5259 -2550 5293
rect -2608 5225 -2596 5259
rect -2562 5225 -2550 5259
rect -2608 5191 -2550 5225
rect -2608 5157 -2596 5191
rect -2562 5157 -2550 5191
rect -2608 5123 -2550 5157
rect -2608 5089 -2596 5123
rect -2562 5089 -2550 5123
rect -2608 5055 -2550 5089
rect -2608 5021 -2596 5055
rect -2562 5021 -2550 5055
rect -2608 4987 -2550 5021
rect -2608 4953 -2596 4987
rect -2562 4953 -2550 4987
rect -2608 4919 -2550 4953
rect -2608 4885 -2596 4919
rect -2562 4885 -2550 4919
rect -2608 4851 -2550 4885
rect -2608 4817 -2596 4851
rect -2562 4817 -2550 4851
rect -2608 4783 -2550 4817
rect -2608 4749 -2596 4783
rect -2562 4749 -2550 4783
rect -2608 4715 -2550 4749
rect -2608 4681 -2596 4715
rect -2562 4681 -2550 4715
rect -2608 4647 -2550 4681
rect -2608 4613 -2596 4647
rect -2562 4613 -2550 4647
rect -2608 4579 -2550 4613
rect -2608 4545 -2596 4579
rect -2562 4545 -2550 4579
rect -2608 4511 -2550 4545
rect -2608 4477 -2596 4511
rect -2562 4477 -2550 4511
rect -2608 4443 -2550 4477
rect -2608 4409 -2596 4443
rect -2562 4409 -2550 4443
rect -2608 4375 -2550 4409
rect -2608 4341 -2596 4375
rect -2562 4341 -2550 4375
rect -2608 4307 -2550 4341
rect -2608 4273 -2596 4307
rect -2562 4273 -2550 4307
rect -2608 4239 -2550 4273
rect -2608 4205 -2596 4239
rect -2562 4205 -2550 4239
rect -2608 4171 -2550 4205
rect -2608 4137 -2596 4171
rect -2562 4137 -2550 4171
rect -2608 4103 -2550 4137
rect -2608 4069 -2596 4103
rect -2562 4069 -2550 4103
rect -2608 4035 -2550 4069
rect -2608 4001 -2596 4035
rect -2562 4001 -2550 4035
rect -2608 3967 -2550 4001
rect -2608 3933 -2596 3967
rect -2562 3933 -2550 3967
rect -2608 3899 -2550 3933
rect -2608 3865 -2596 3899
rect -2562 3865 -2550 3899
rect -2608 3831 -2550 3865
rect -2608 3797 -2596 3831
rect -2562 3797 -2550 3831
rect -2608 3763 -2550 3797
rect -2608 3729 -2596 3763
rect -2562 3729 -2550 3763
rect -2608 3695 -2550 3729
rect -2608 3661 -2596 3695
rect -2562 3661 -2550 3695
rect -2608 3630 -2550 3661
rect -2166 5599 -2108 5630
rect -2166 5565 -2154 5599
rect -2120 5565 -2108 5599
rect -2166 5531 -2108 5565
rect -2166 5497 -2154 5531
rect -2120 5497 -2108 5531
rect -2166 5463 -2108 5497
rect -2166 5429 -2154 5463
rect -2120 5429 -2108 5463
rect -2166 5395 -2108 5429
rect -2166 5361 -2154 5395
rect -2120 5361 -2108 5395
rect -2166 5327 -2108 5361
rect -2166 5293 -2154 5327
rect -2120 5293 -2108 5327
rect -2166 5259 -2108 5293
rect -2166 5225 -2154 5259
rect -2120 5225 -2108 5259
rect -2166 5191 -2108 5225
rect -2166 5157 -2154 5191
rect -2120 5157 -2108 5191
rect -2166 5123 -2108 5157
rect -2166 5089 -2154 5123
rect -2120 5089 -2108 5123
rect -2166 5055 -2108 5089
rect -2166 5021 -2154 5055
rect -2120 5021 -2108 5055
rect -2166 4987 -2108 5021
rect -2166 4953 -2154 4987
rect -2120 4953 -2108 4987
rect -2166 4919 -2108 4953
rect -2166 4885 -2154 4919
rect -2120 4885 -2108 4919
rect -2166 4851 -2108 4885
rect -2166 4817 -2154 4851
rect -2120 4817 -2108 4851
rect -2166 4783 -2108 4817
rect -2166 4749 -2154 4783
rect -2120 4749 -2108 4783
rect -2166 4715 -2108 4749
rect -2166 4681 -2154 4715
rect -2120 4681 -2108 4715
rect -2166 4647 -2108 4681
rect -2166 4613 -2154 4647
rect -2120 4613 -2108 4647
rect -2166 4579 -2108 4613
rect -2166 4545 -2154 4579
rect -2120 4545 -2108 4579
rect -2166 4511 -2108 4545
rect -2166 4477 -2154 4511
rect -2120 4477 -2108 4511
rect -2166 4443 -2108 4477
rect -2166 4409 -2154 4443
rect -2120 4409 -2108 4443
rect -2166 4375 -2108 4409
rect -2166 4341 -2154 4375
rect -2120 4341 -2108 4375
rect -2166 4307 -2108 4341
rect -2166 4273 -2154 4307
rect -2120 4273 -2108 4307
rect -2166 4239 -2108 4273
rect -2166 4205 -2154 4239
rect -2120 4205 -2108 4239
rect -2166 4171 -2108 4205
rect -2166 4137 -2154 4171
rect -2120 4137 -2108 4171
rect -2166 4103 -2108 4137
rect -2166 4069 -2154 4103
rect -2120 4069 -2108 4103
rect -2166 4035 -2108 4069
rect -2166 4001 -2154 4035
rect -2120 4001 -2108 4035
rect -2166 3967 -2108 4001
rect -2166 3933 -2154 3967
rect -2120 3933 -2108 3967
rect -2166 3899 -2108 3933
rect -2166 3865 -2154 3899
rect -2120 3865 -2108 3899
rect -2166 3831 -2108 3865
rect -2166 3797 -2154 3831
rect -2120 3797 -2108 3831
rect -2166 3763 -2108 3797
rect -2166 3729 -2154 3763
rect -2120 3729 -2108 3763
rect -2166 3695 -2108 3729
rect -2166 3661 -2154 3695
rect -2120 3661 -2108 3695
rect -2166 3630 -2108 3661
rect -1908 5599 -1850 5630
rect -1908 5565 -1896 5599
rect -1862 5565 -1850 5599
rect -1908 5531 -1850 5565
rect -1908 5497 -1896 5531
rect -1862 5497 -1850 5531
rect -1908 5463 -1850 5497
rect -1908 5429 -1896 5463
rect -1862 5429 -1850 5463
rect -1908 5395 -1850 5429
rect -1908 5361 -1896 5395
rect -1862 5361 -1850 5395
rect -1908 5327 -1850 5361
rect -1908 5293 -1896 5327
rect -1862 5293 -1850 5327
rect -1908 5259 -1850 5293
rect -1908 5225 -1896 5259
rect -1862 5225 -1850 5259
rect -1908 5191 -1850 5225
rect -1908 5157 -1896 5191
rect -1862 5157 -1850 5191
rect -1908 5123 -1850 5157
rect -1908 5089 -1896 5123
rect -1862 5089 -1850 5123
rect -1908 5055 -1850 5089
rect -1908 5021 -1896 5055
rect -1862 5021 -1850 5055
rect -1908 4987 -1850 5021
rect -1908 4953 -1896 4987
rect -1862 4953 -1850 4987
rect -1908 4919 -1850 4953
rect -1908 4885 -1896 4919
rect -1862 4885 -1850 4919
rect -1908 4851 -1850 4885
rect -1908 4817 -1896 4851
rect -1862 4817 -1850 4851
rect -1908 4783 -1850 4817
rect -1908 4749 -1896 4783
rect -1862 4749 -1850 4783
rect -1908 4715 -1850 4749
rect -1908 4681 -1896 4715
rect -1862 4681 -1850 4715
rect -1908 4647 -1850 4681
rect -1908 4613 -1896 4647
rect -1862 4613 -1850 4647
rect -1908 4579 -1850 4613
rect -1908 4545 -1896 4579
rect -1862 4545 -1850 4579
rect -1908 4511 -1850 4545
rect -1908 4477 -1896 4511
rect -1862 4477 -1850 4511
rect -1908 4443 -1850 4477
rect -1908 4409 -1896 4443
rect -1862 4409 -1850 4443
rect -1908 4375 -1850 4409
rect -1908 4341 -1896 4375
rect -1862 4341 -1850 4375
rect -1908 4307 -1850 4341
rect -1908 4273 -1896 4307
rect -1862 4273 -1850 4307
rect -1908 4239 -1850 4273
rect -1908 4205 -1896 4239
rect -1862 4205 -1850 4239
rect -1908 4171 -1850 4205
rect -1908 4137 -1896 4171
rect -1862 4137 -1850 4171
rect -1908 4103 -1850 4137
rect -1908 4069 -1896 4103
rect -1862 4069 -1850 4103
rect -1908 4035 -1850 4069
rect -1908 4001 -1896 4035
rect -1862 4001 -1850 4035
rect -1908 3967 -1850 4001
rect -1908 3933 -1896 3967
rect -1862 3933 -1850 3967
rect -1908 3899 -1850 3933
rect -1908 3865 -1896 3899
rect -1862 3865 -1850 3899
rect -1908 3831 -1850 3865
rect -1908 3797 -1896 3831
rect -1862 3797 -1850 3831
rect -1908 3763 -1850 3797
rect -1908 3729 -1896 3763
rect -1862 3729 -1850 3763
rect -1908 3695 -1850 3729
rect -1908 3661 -1896 3695
rect -1862 3661 -1850 3695
rect -1908 3630 -1850 3661
rect -1466 5599 -1408 5630
rect -1466 5565 -1454 5599
rect -1420 5565 -1408 5599
rect -1466 5531 -1408 5565
rect -1466 5497 -1454 5531
rect -1420 5497 -1408 5531
rect -1466 5463 -1408 5497
rect -1466 5429 -1454 5463
rect -1420 5429 -1408 5463
rect -1466 5395 -1408 5429
rect -1466 5361 -1454 5395
rect -1420 5361 -1408 5395
rect -1466 5327 -1408 5361
rect -1466 5293 -1454 5327
rect -1420 5293 -1408 5327
rect -1466 5259 -1408 5293
rect -1466 5225 -1454 5259
rect -1420 5225 -1408 5259
rect -1466 5191 -1408 5225
rect -1466 5157 -1454 5191
rect -1420 5157 -1408 5191
rect -1466 5123 -1408 5157
rect -1466 5089 -1454 5123
rect -1420 5089 -1408 5123
rect -1466 5055 -1408 5089
rect -1466 5021 -1454 5055
rect -1420 5021 -1408 5055
rect -1466 4987 -1408 5021
rect -1466 4953 -1454 4987
rect -1420 4953 -1408 4987
rect -1466 4919 -1408 4953
rect -1466 4885 -1454 4919
rect -1420 4885 -1408 4919
rect -1466 4851 -1408 4885
rect -1466 4817 -1454 4851
rect -1420 4817 -1408 4851
rect -1466 4783 -1408 4817
rect -1466 4749 -1454 4783
rect -1420 4749 -1408 4783
rect -1466 4715 -1408 4749
rect -1466 4681 -1454 4715
rect -1420 4681 -1408 4715
rect -1466 4647 -1408 4681
rect -1466 4613 -1454 4647
rect -1420 4613 -1408 4647
rect -1466 4579 -1408 4613
rect -1466 4545 -1454 4579
rect -1420 4545 -1408 4579
rect -1466 4511 -1408 4545
rect -1466 4477 -1454 4511
rect -1420 4477 -1408 4511
rect -1466 4443 -1408 4477
rect -1466 4409 -1454 4443
rect -1420 4409 -1408 4443
rect -1466 4375 -1408 4409
rect -1466 4341 -1454 4375
rect -1420 4341 -1408 4375
rect -1466 4307 -1408 4341
rect -1466 4273 -1454 4307
rect -1420 4273 -1408 4307
rect -1466 4239 -1408 4273
rect -1466 4205 -1454 4239
rect -1420 4205 -1408 4239
rect -1466 4171 -1408 4205
rect -1466 4137 -1454 4171
rect -1420 4137 -1408 4171
rect -1466 4103 -1408 4137
rect -1466 4069 -1454 4103
rect -1420 4069 -1408 4103
rect -1466 4035 -1408 4069
rect -1466 4001 -1454 4035
rect -1420 4001 -1408 4035
rect -1466 3967 -1408 4001
rect -1466 3933 -1454 3967
rect -1420 3933 -1408 3967
rect -1466 3899 -1408 3933
rect -1466 3865 -1454 3899
rect -1420 3865 -1408 3899
rect -1466 3831 -1408 3865
rect -1466 3797 -1454 3831
rect -1420 3797 -1408 3831
rect -1466 3763 -1408 3797
rect -1466 3729 -1454 3763
rect -1420 3729 -1408 3763
rect -1466 3695 -1408 3729
rect -1466 3661 -1454 3695
rect -1420 3661 -1408 3695
rect -1466 3630 -1408 3661
rect -1208 5599 -1150 5630
rect -1208 5565 -1196 5599
rect -1162 5565 -1150 5599
rect -1208 5531 -1150 5565
rect -1208 5497 -1196 5531
rect -1162 5497 -1150 5531
rect -1208 5463 -1150 5497
rect -1208 5429 -1196 5463
rect -1162 5429 -1150 5463
rect -1208 5395 -1150 5429
rect -1208 5361 -1196 5395
rect -1162 5361 -1150 5395
rect -1208 5327 -1150 5361
rect -1208 5293 -1196 5327
rect -1162 5293 -1150 5327
rect -1208 5259 -1150 5293
rect -1208 5225 -1196 5259
rect -1162 5225 -1150 5259
rect -1208 5191 -1150 5225
rect -1208 5157 -1196 5191
rect -1162 5157 -1150 5191
rect -1208 5123 -1150 5157
rect -1208 5089 -1196 5123
rect -1162 5089 -1150 5123
rect -1208 5055 -1150 5089
rect -1208 5021 -1196 5055
rect -1162 5021 -1150 5055
rect -1208 4987 -1150 5021
rect -1208 4953 -1196 4987
rect -1162 4953 -1150 4987
rect -1208 4919 -1150 4953
rect -1208 4885 -1196 4919
rect -1162 4885 -1150 4919
rect -1208 4851 -1150 4885
rect -1208 4817 -1196 4851
rect -1162 4817 -1150 4851
rect -1208 4783 -1150 4817
rect -1208 4749 -1196 4783
rect -1162 4749 -1150 4783
rect -1208 4715 -1150 4749
rect -1208 4681 -1196 4715
rect -1162 4681 -1150 4715
rect -1208 4647 -1150 4681
rect -1208 4613 -1196 4647
rect -1162 4613 -1150 4647
rect -1208 4579 -1150 4613
rect -1208 4545 -1196 4579
rect -1162 4545 -1150 4579
rect -1208 4511 -1150 4545
rect -1208 4477 -1196 4511
rect -1162 4477 -1150 4511
rect -1208 4443 -1150 4477
rect -1208 4409 -1196 4443
rect -1162 4409 -1150 4443
rect -1208 4375 -1150 4409
rect -1208 4341 -1196 4375
rect -1162 4341 -1150 4375
rect -1208 4307 -1150 4341
rect -1208 4273 -1196 4307
rect -1162 4273 -1150 4307
rect -1208 4239 -1150 4273
rect -1208 4205 -1196 4239
rect -1162 4205 -1150 4239
rect -1208 4171 -1150 4205
rect -1208 4137 -1196 4171
rect -1162 4137 -1150 4171
rect -1208 4103 -1150 4137
rect -1208 4069 -1196 4103
rect -1162 4069 -1150 4103
rect -1208 4035 -1150 4069
rect -1208 4001 -1196 4035
rect -1162 4001 -1150 4035
rect -1208 3967 -1150 4001
rect -1208 3933 -1196 3967
rect -1162 3933 -1150 3967
rect -1208 3899 -1150 3933
rect -1208 3865 -1196 3899
rect -1162 3865 -1150 3899
rect -1208 3831 -1150 3865
rect -1208 3797 -1196 3831
rect -1162 3797 -1150 3831
rect -1208 3763 -1150 3797
rect -1208 3729 -1196 3763
rect -1162 3729 -1150 3763
rect -1208 3695 -1150 3729
rect -1208 3661 -1196 3695
rect -1162 3661 -1150 3695
rect -1208 3630 -1150 3661
rect -766 5599 -708 5630
rect -766 5565 -754 5599
rect -720 5565 -708 5599
rect -766 5531 -708 5565
rect -766 5497 -754 5531
rect -720 5497 -708 5531
rect -766 5463 -708 5497
rect -766 5429 -754 5463
rect -720 5429 -708 5463
rect -766 5395 -708 5429
rect -766 5361 -754 5395
rect -720 5361 -708 5395
rect -766 5327 -708 5361
rect -766 5293 -754 5327
rect -720 5293 -708 5327
rect -766 5259 -708 5293
rect -766 5225 -754 5259
rect -720 5225 -708 5259
rect -766 5191 -708 5225
rect -766 5157 -754 5191
rect -720 5157 -708 5191
rect -766 5123 -708 5157
rect -766 5089 -754 5123
rect -720 5089 -708 5123
rect -766 5055 -708 5089
rect -766 5021 -754 5055
rect -720 5021 -708 5055
rect -766 4987 -708 5021
rect -766 4953 -754 4987
rect -720 4953 -708 4987
rect -766 4919 -708 4953
rect -766 4885 -754 4919
rect -720 4885 -708 4919
rect -766 4851 -708 4885
rect -766 4817 -754 4851
rect -720 4817 -708 4851
rect -766 4783 -708 4817
rect -766 4749 -754 4783
rect -720 4749 -708 4783
rect -766 4715 -708 4749
rect -766 4681 -754 4715
rect -720 4681 -708 4715
rect -766 4647 -708 4681
rect -766 4613 -754 4647
rect -720 4613 -708 4647
rect -766 4579 -708 4613
rect -766 4545 -754 4579
rect -720 4545 -708 4579
rect -766 4511 -708 4545
rect -766 4477 -754 4511
rect -720 4477 -708 4511
rect -766 4443 -708 4477
rect -766 4409 -754 4443
rect -720 4409 -708 4443
rect -766 4375 -708 4409
rect -766 4341 -754 4375
rect -720 4341 -708 4375
rect -766 4307 -708 4341
rect -766 4273 -754 4307
rect -720 4273 -708 4307
rect -766 4239 -708 4273
rect -766 4205 -754 4239
rect -720 4205 -708 4239
rect -766 4171 -708 4205
rect -766 4137 -754 4171
rect -720 4137 -708 4171
rect -766 4103 -708 4137
rect -766 4069 -754 4103
rect -720 4069 -708 4103
rect -766 4035 -708 4069
rect -766 4001 -754 4035
rect -720 4001 -708 4035
rect -766 3967 -708 4001
rect -766 3933 -754 3967
rect -720 3933 -708 3967
rect -766 3899 -708 3933
rect -766 3865 -754 3899
rect -720 3865 -708 3899
rect -766 3831 -708 3865
rect -766 3797 -754 3831
rect -720 3797 -708 3831
rect -766 3763 -708 3797
rect -766 3729 -754 3763
rect -720 3729 -708 3763
rect -766 3695 -708 3729
rect -766 3661 -754 3695
rect -720 3661 -708 3695
rect -766 3630 -708 3661
rect -508 5599 -450 5630
rect -508 5565 -496 5599
rect -462 5565 -450 5599
rect -508 5531 -450 5565
rect -508 5497 -496 5531
rect -462 5497 -450 5531
rect -508 5463 -450 5497
rect -508 5429 -496 5463
rect -462 5429 -450 5463
rect -508 5395 -450 5429
rect -508 5361 -496 5395
rect -462 5361 -450 5395
rect -508 5327 -450 5361
rect -508 5293 -496 5327
rect -462 5293 -450 5327
rect -508 5259 -450 5293
rect -508 5225 -496 5259
rect -462 5225 -450 5259
rect -508 5191 -450 5225
rect -508 5157 -496 5191
rect -462 5157 -450 5191
rect -508 5123 -450 5157
rect -508 5089 -496 5123
rect -462 5089 -450 5123
rect -508 5055 -450 5089
rect -508 5021 -496 5055
rect -462 5021 -450 5055
rect -508 4987 -450 5021
rect -508 4953 -496 4987
rect -462 4953 -450 4987
rect -508 4919 -450 4953
rect -508 4885 -496 4919
rect -462 4885 -450 4919
rect -508 4851 -450 4885
rect -508 4817 -496 4851
rect -462 4817 -450 4851
rect -508 4783 -450 4817
rect -508 4749 -496 4783
rect -462 4749 -450 4783
rect -508 4715 -450 4749
rect -508 4681 -496 4715
rect -462 4681 -450 4715
rect -508 4647 -450 4681
rect -508 4613 -496 4647
rect -462 4613 -450 4647
rect -508 4579 -450 4613
rect -508 4545 -496 4579
rect -462 4545 -450 4579
rect -508 4511 -450 4545
rect -508 4477 -496 4511
rect -462 4477 -450 4511
rect -508 4443 -450 4477
rect -508 4409 -496 4443
rect -462 4409 -450 4443
rect -508 4375 -450 4409
rect -508 4341 -496 4375
rect -462 4341 -450 4375
rect -508 4307 -450 4341
rect -508 4273 -496 4307
rect -462 4273 -450 4307
rect -508 4239 -450 4273
rect -508 4205 -496 4239
rect -462 4205 -450 4239
rect -508 4171 -450 4205
rect -508 4137 -496 4171
rect -462 4137 -450 4171
rect -508 4103 -450 4137
rect -508 4069 -496 4103
rect -462 4069 -450 4103
rect -508 4035 -450 4069
rect -508 4001 -496 4035
rect -462 4001 -450 4035
rect -508 3967 -450 4001
rect -508 3933 -496 3967
rect -462 3933 -450 3967
rect -508 3899 -450 3933
rect -508 3865 -496 3899
rect -462 3865 -450 3899
rect -508 3831 -450 3865
rect -508 3797 -496 3831
rect -462 3797 -450 3831
rect -508 3763 -450 3797
rect -508 3729 -496 3763
rect -462 3729 -450 3763
rect -508 3695 -450 3729
rect -508 3661 -496 3695
rect -462 3661 -450 3695
rect -508 3630 -450 3661
rect -66 5599 -8 5630
rect -66 5565 -54 5599
rect -20 5565 -8 5599
rect -66 5531 -8 5565
rect -66 5497 -54 5531
rect -20 5497 -8 5531
rect -66 5463 -8 5497
rect -66 5429 -54 5463
rect -20 5429 -8 5463
rect -66 5395 -8 5429
rect -66 5361 -54 5395
rect -20 5361 -8 5395
rect -66 5327 -8 5361
rect -66 5293 -54 5327
rect -20 5293 -8 5327
rect -66 5259 -8 5293
rect -66 5225 -54 5259
rect -20 5225 -8 5259
rect -66 5191 -8 5225
rect -66 5157 -54 5191
rect -20 5157 -8 5191
rect -66 5123 -8 5157
rect -66 5089 -54 5123
rect -20 5089 -8 5123
rect -66 5055 -8 5089
rect -66 5021 -54 5055
rect -20 5021 -8 5055
rect -66 4987 -8 5021
rect -66 4953 -54 4987
rect -20 4953 -8 4987
rect -66 4919 -8 4953
rect -66 4885 -54 4919
rect -20 4885 -8 4919
rect -66 4851 -8 4885
rect -66 4817 -54 4851
rect -20 4817 -8 4851
rect -66 4783 -8 4817
rect -66 4749 -54 4783
rect -20 4749 -8 4783
rect -66 4715 -8 4749
rect -66 4681 -54 4715
rect -20 4681 -8 4715
rect -66 4647 -8 4681
rect -66 4613 -54 4647
rect -20 4613 -8 4647
rect -66 4579 -8 4613
rect -66 4545 -54 4579
rect -20 4545 -8 4579
rect -66 4511 -8 4545
rect -66 4477 -54 4511
rect -20 4477 -8 4511
rect -66 4443 -8 4477
rect -66 4409 -54 4443
rect -20 4409 -8 4443
rect -66 4375 -8 4409
rect -66 4341 -54 4375
rect -20 4341 -8 4375
rect -66 4307 -8 4341
rect -66 4273 -54 4307
rect -20 4273 -8 4307
rect -66 4239 -8 4273
rect -66 4205 -54 4239
rect -20 4205 -8 4239
rect -66 4171 -8 4205
rect -66 4137 -54 4171
rect -20 4137 -8 4171
rect -66 4103 -8 4137
rect -66 4069 -54 4103
rect -20 4069 -8 4103
rect -66 4035 -8 4069
rect -66 4001 -54 4035
rect -20 4001 -8 4035
rect -66 3967 -8 4001
rect -66 3933 -54 3967
rect -20 3933 -8 3967
rect -66 3899 -8 3933
rect -66 3865 -54 3899
rect -20 3865 -8 3899
rect -66 3831 -8 3865
rect -66 3797 -54 3831
rect -20 3797 -8 3831
rect -66 3763 -8 3797
rect -66 3729 -54 3763
rect -20 3729 -8 3763
rect -66 3695 -8 3729
rect -66 3661 -54 3695
rect -20 3661 -8 3695
rect -66 3630 -8 3661
rect 192 5599 250 5630
rect 192 5565 204 5599
rect 238 5565 250 5599
rect 192 5531 250 5565
rect 192 5497 204 5531
rect 238 5497 250 5531
rect 192 5463 250 5497
rect 192 5429 204 5463
rect 238 5429 250 5463
rect 192 5395 250 5429
rect 192 5361 204 5395
rect 238 5361 250 5395
rect 192 5327 250 5361
rect 192 5293 204 5327
rect 238 5293 250 5327
rect 192 5259 250 5293
rect 192 5225 204 5259
rect 238 5225 250 5259
rect 192 5191 250 5225
rect 192 5157 204 5191
rect 238 5157 250 5191
rect 192 5123 250 5157
rect 192 5089 204 5123
rect 238 5089 250 5123
rect 192 5055 250 5089
rect 192 5021 204 5055
rect 238 5021 250 5055
rect 192 4987 250 5021
rect 192 4953 204 4987
rect 238 4953 250 4987
rect 192 4919 250 4953
rect 192 4885 204 4919
rect 238 4885 250 4919
rect 192 4851 250 4885
rect 192 4817 204 4851
rect 238 4817 250 4851
rect 192 4783 250 4817
rect 192 4749 204 4783
rect 238 4749 250 4783
rect 192 4715 250 4749
rect 192 4681 204 4715
rect 238 4681 250 4715
rect 192 4647 250 4681
rect 192 4613 204 4647
rect 238 4613 250 4647
rect 192 4579 250 4613
rect 192 4545 204 4579
rect 238 4545 250 4579
rect 192 4511 250 4545
rect 192 4477 204 4511
rect 238 4477 250 4511
rect 192 4443 250 4477
rect 192 4409 204 4443
rect 238 4409 250 4443
rect 192 4375 250 4409
rect 192 4341 204 4375
rect 238 4341 250 4375
rect 192 4307 250 4341
rect 192 4273 204 4307
rect 238 4273 250 4307
rect 192 4239 250 4273
rect 192 4205 204 4239
rect 238 4205 250 4239
rect 192 4171 250 4205
rect 192 4137 204 4171
rect 238 4137 250 4171
rect 192 4103 250 4137
rect 192 4069 204 4103
rect 238 4069 250 4103
rect 192 4035 250 4069
rect 192 4001 204 4035
rect 238 4001 250 4035
rect 192 3967 250 4001
rect 192 3933 204 3967
rect 238 3933 250 3967
rect 192 3899 250 3933
rect 192 3865 204 3899
rect 238 3865 250 3899
rect 192 3831 250 3865
rect 192 3797 204 3831
rect 238 3797 250 3831
rect 192 3763 250 3797
rect 192 3729 204 3763
rect 238 3729 250 3763
rect 192 3695 250 3729
rect 192 3661 204 3695
rect 238 3661 250 3695
rect 192 3630 250 3661
rect 634 5599 692 5630
rect 634 5565 646 5599
rect 680 5565 692 5599
rect 634 5531 692 5565
rect 634 5497 646 5531
rect 680 5497 692 5531
rect 634 5463 692 5497
rect 634 5429 646 5463
rect 680 5429 692 5463
rect 634 5395 692 5429
rect 634 5361 646 5395
rect 680 5361 692 5395
rect 634 5327 692 5361
rect 634 5293 646 5327
rect 680 5293 692 5327
rect 634 5259 692 5293
rect 634 5225 646 5259
rect 680 5225 692 5259
rect 634 5191 692 5225
rect 634 5157 646 5191
rect 680 5157 692 5191
rect 634 5123 692 5157
rect 634 5089 646 5123
rect 680 5089 692 5123
rect 634 5055 692 5089
rect 634 5021 646 5055
rect 680 5021 692 5055
rect 634 4987 692 5021
rect 634 4953 646 4987
rect 680 4953 692 4987
rect 634 4919 692 4953
rect 634 4885 646 4919
rect 680 4885 692 4919
rect 634 4851 692 4885
rect 634 4817 646 4851
rect 680 4817 692 4851
rect 634 4783 692 4817
rect 634 4749 646 4783
rect 680 4749 692 4783
rect 634 4715 692 4749
rect 634 4681 646 4715
rect 680 4681 692 4715
rect 634 4647 692 4681
rect 634 4613 646 4647
rect 680 4613 692 4647
rect 634 4579 692 4613
rect 634 4545 646 4579
rect 680 4545 692 4579
rect 634 4511 692 4545
rect 634 4477 646 4511
rect 680 4477 692 4511
rect 634 4443 692 4477
rect 634 4409 646 4443
rect 680 4409 692 4443
rect 634 4375 692 4409
rect 634 4341 646 4375
rect 680 4341 692 4375
rect 634 4307 692 4341
rect 634 4273 646 4307
rect 680 4273 692 4307
rect 634 4239 692 4273
rect 634 4205 646 4239
rect 680 4205 692 4239
rect 634 4171 692 4205
rect 634 4137 646 4171
rect 680 4137 692 4171
rect 634 4103 692 4137
rect 634 4069 646 4103
rect 680 4069 692 4103
rect 634 4035 692 4069
rect 634 4001 646 4035
rect 680 4001 692 4035
rect 634 3967 692 4001
rect 634 3933 646 3967
rect 680 3933 692 3967
rect 634 3899 692 3933
rect 634 3865 646 3899
rect 680 3865 692 3899
rect 634 3831 692 3865
rect 634 3797 646 3831
rect 680 3797 692 3831
rect 634 3763 692 3797
rect 634 3729 646 3763
rect 680 3729 692 3763
rect 634 3695 692 3729
rect 634 3661 646 3695
rect 680 3661 692 3695
rect 634 3630 692 3661
rect 892 5599 950 5630
rect 892 5565 904 5599
rect 938 5565 950 5599
rect 892 5531 950 5565
rect 892 5497 904 5531
rect 938 5497 950 5531
rect 892 5463 950 5497
rect 892 5429 904 5463
rect 938 5429 950 5463
rect 892 5395 950 5429
rect 892 5361 904 5395
rect 938 5361 950 5395
rect 892 5327 950 5361
rect 892 5293 904 5327
rect 938 5293 950 5327
rect 892 5259 950 5293
rect 892 5225 904 5259
rect 938 5225 950 5259
rect 892 5191 950 5225
rect 892 5157 904 5191
rect 938 5157 950 5191
rect 892 5123 950 5157
rect 892 5089 904 5123
rect 938 5089 950 5123
rect 892 5055 950 5089
rect 892 5021 904 5055
rect 938 5021 950 5055
rect 892 4987 950 5021
rect 892 4953 904 4987
rect 938 4953 950 4987
rect 892 4919 950 4953
rect 892 4885 904 4919
rect 938 4885 950 4919
rect 892 4851 950 4885
rect 892 4817 904 4851
rect 938 4817 950 4851
rect 892 4783 950 4817
rect 892 4749 904 4783
rect 938 4749 950 4783
rect 892 4715 950 4749
rect 892 4681 904 4715
rect 938 4681 950 4715
rect 892 4647 950 4681
rect 892 4613 904 4647
rect 938 4613 950 4647
rect 892 4579 950 4613
rect 892 4545 904 4579
rect 938 4545 950 4579
rect 892 4511 950 4545
rect 892 4477 904 4511
rect 938 4477 950 4511
rect 892 4443 950 4477
rect 892 4409 904 4443
rect 938 4409 950 4443
rect 892 4375 950 4409
rect 892 4341 904 4375
rect 938 4341 950 4375
rect 892 4307 950 4341
rect 892 4273 904 4307
rect 938 4273 950 4307
rect 892 4239 950 4273
rect 892 4205 904 4239
rect 938 4205 950 4239
rect 892 4171 950 4205
rect 892 4137 904 4171
rect 938 4137 950 4171
rect 892 4103 950 4137
rect 892 4069 904 4103
rect 938 4069 950 4103
rect 892 4035 950 4069
rect 892 4001 904 4035
rect 938 4001 950 4035
rect 892 3967 950 4001
rect 892 3933 904 3967
rect 938 3933 950 3967
rect 892 3899 950 3933
rect 892 3865 904 3899
rect 938 3865 950 3899
rect 892 3831 950 3865
rect 892 3797 904 3831
rect 938 3797 950 3831
rect 892 3763 950 3797
rect 892 3729 904 3763
rect 938 3729 950 3763
rect 892 3695 950 3729
rect 892 3661 904 3695
rect 938 3661 950 3695
rect 892 3630 950 3661
rect 1334 5599 1392 5630
rect 1334 5565 1346 5599
rect 1380 5565 1392 5599
rect 1334 5531 1392 5565
rect 1334 5497 1346 5531
rect 1380 5497 1392 5531
rect 1334 5463 1392 5497
rect 1334 5429 1346 5463
rect 1380 5429 1392 5463
rect 1334 5395 1392 5429
rect 1334 5361 1346 5395
rect 1380 5361 1392 5395
rect 1334 5327 1392 5361
rect 1334 5293 1346 5327
rect 1380 5293 1392 5327
rect 1334 5259 1392 5293
rect 1334 5225 1346 5259
rect 1380 5225 1392 5259
rect 1334 5191 1392 5225
rect 1334 5157 1346 5191
rect 1380 5157 1392 5191
rect 1334 5123 1392 5157
rect 1334 5089 1346 5123
rect 1380 5089 1392 5123
rect 1334 5055 1392 5089
rect 1334 5021 1346 5055
rect 1380 5021 1392 5055
rect 1334 4987 1392 5021
rect 1334 4953 1346 4987
rect 1380 4953 1392 4987
rect 1334 4919 1392 4953
rect 1334 4885 1346 4919
rect 1380 4885 1392 4919
rect 1334 4851 1392 4885
rect 1334 4817 1346 4851
rect 1380 4817 1392 4851
rect 1334 4783 1392 4817
rect 1334 4749 1346 4783
rect 1380 4749 1392 4783
rect 1334 4715 1392 4749
rect 1334 4681 1346 4715
rect 1380 4681 1392 4715
rect 1334 4647 1392 4681
rect 1334 4613 1346 4647
rect 1380 4613 1392 4647
rect 1334 4579 1392 4613
rect 1334 4545 1346 4579
rect 1380 4545 1392 4579
rect 1334 4511 1392 4545
rect 1334 4477 1346 4511
rect 1380 4477 1392 4511
rect 1334 4443 1392 4477
rect 1334 4409 1346 4443
rect 1380 4409 1392 4443
rect 1334 4375 1392 4409
rect 1334 4341 1346 4375
rect 1380 4341 1392 4375
rect 1334 4307 1392 4341
rect 1334 4273 1346 4307
rect 1380 4273 1392 4307
rect 1334 4239 1392 4273
rect 1334 4205 1346 4239
rect 1380 4205 1392 4239
rect 1334 4171 1392 4205
rect 1334 4137 1346 4171
rect 1380 4137 1392 4171
rect 1334 4103 1392 4137
rect 1334 4069 1346 4103
rect 1380 4069 1392 4103
rect 1334 4035 1392 4069
rect 1334 4001 1346 4035
rect 1380 4001 1392 4035
rect 1334 3967 1392 4001
rect 1334 3933 1346 3967
rect 1380 3933 1392 3967
rect 1334 3899 1392 3933
rect 1334 3865 1346 3899
rect 1380 3865 1392 3899
rect 1334 3831 1392 3865
rect 1334 3797 1346 3831
rect 1380 3797 1392 3831
rect 1334 3763 1392 3797
rect 1334 3729 1346 3763
rect 1380 3729 1392 3763
rect 1334 3695 1392 3729
rect 1334 3661 1346 3695
rect 1380 3661 1392 3695
rect 1334 3630 1392 3661
rect 1592 5599 1650 5630
rect 1592 5565 1604 5599
rect 1638 5565 1650 5599
rect 1592 5531 1650 5565
rect 1592 5497 1604 5531
rect 1638 5497 1650 5531
rect 1592 5463 1650 5497
rect 1592 5429 1604 5463
rect 1638 5429 1650 5463
rect 1592 5395 1650 5429
rect 1592 5361 1604 5395
rect 1638 5361 1650 5395
rect 1592 5327 1650 5361
rect 1592 5293 1604 5327
rect 1638 5293 1650 5327
rect 1592 5259 1650 5293
rect 1592 5225 1604 5259
rect 1638 5225 1650 5259
rect 1592 5191 1650 5225
rect 1592 5157 1604 5191
rect 1638 5157 1650 5191
rect 1592 5123 1650 5157
rect 1592 5089 1604 5123
rect 1638 5089 1650 5123
rect 1592 5055 1650 5089
rect 1592 5021 1604 5055
rect 1638 5021 1650 5055
rect 1592 4987 1650 5021
rect 1592 4953 1604 4987
rect 1638 4953 1650 4987
rect 1592 4919 1650 4953
rect 1592 4885 1604 4919
rect 1638 4885 1650 4919
rect 1592 4851 1650 4885
rect 1592 4817 1604 4851
rect 1638 4817 1650 4851
rect 1592 4783 1650 4817
rect 1592 4749 1604 4783
rect 1638 4749 1650 4783
rect 1592 4715 1650 4749
rect 1592 4681 1604 4715
rect 1638 4681 1650 4715
rect 1592 4647 1650 4681
rect 1592 4613 1604 4647
rect 1638 4613 1650 4647
rect 1592 4579 1650 4613
rect 1592 4545 1604 4579
rect 1638 4545 1650 4579
rect 1592 4511 1650 4545
rect 1592 4477 1604 4511
rect 1638 4477 1650 4511
rect 1592 4443 1650 4477
rect 1592 4409 1604 4443
rect 1638 4409 1650 4443
rect 1592 4375 1650 4409
rect 1592 4341 1604 4375
rect 1638 4341 1650 4375
rect 1592 4307 1650 4341
rect 1592 4273 1604 4307
rect 1638 4273 1650 4307
rect 1592 4239 1650 4273
rect 1592 4205 1604 4239
rect 1638 4205 1650 4239
rect 1592 4171 1650 4205
rect 1592 4137 1604 4171
rect 1638 4137 1650 4171
rect 1592 4103 1650 4137
rect 1592 4069 1604 4103
rect 1638 4069 1650 4103
rect 1592 4035 1650 4069
rect 1592 4001 1604 4035
rect 1638 4001 1650 4035
rect 1592 3967 1650 4001
rect 1592 3933 1604 3967
rect 1638 3933 1650 3967
rect 1592 3899 1650 3933
rect 1592 3865 1604 3899
rect 1638 3865 1650 3899
rect 1592 3831 1650 3865
rect 1592 3797 1604 3831
rect 1638 3797 1650 3831
rect 1592 3763 1650 3797
rect 1592 3729 1604 3763
rect 1638 3729 1650 3763
rect 1592 3695 1650 3729
rect 1592 3661 1604 3695
rect 1638 3661 1650 3695
rect 1592 3630 1650 3661
rect 2034 5599 2092 5630
rect 2034 5565 2046 5599
rect 2080 5565 2092 5599
rect 2034 5531 2092 5565
rect 2034 5497 2046 5531
rect 2080 5497 2092 5531
rect 2034 5463 2092 5497
rect 2034 5429 2046 5463
rect 2080 5429 2092 5463
rect 2034 5395 2092 5429
rect 2034 5361 2046 5395
rect 2080 5361 2092 5395
rect 2034 5327 2092 5361
rect 2034 5293 2046 5327
rect 2080 5293 2092 5327
rect 2034 5259 2092 5293
rect 2034 5225 2046 5259
rect 2080 5225 2092 5259
rect 2034 5191 2092 5225
rect 2034 5157 2046 5191
rect 2080 5157 2092 5191
rect 2034 5123 2092 5157
rect 2034 5089 2046 5123
rect 2080 5089 2092 5123
rect 2034 5055 2092 5089
rect 2034 5021 2046 5055
rect 2080 5021 2092 5055
rect 2034 4987 2092 5021
rect 2034 4953 2046 4987
rect 2080 4953 2092 4987
rect 2034 4919 2092 4953
rect 2034 4885 2046 4919
rect 2080 4885 2092 4919
rect 2034 4851 2092 4885
rect 2034 4817 2046 4851
rect 2080 4817 2092 4851
rect 2034 4783 2092 4817
rect 2034 4749 2046 4783
rect 2080 4749 2092 4783
rect 2034 4715 2092 4749
rect 2034 4681 2046 4715
rect 2080 4681 2092 4715
rect 2034 4647 2092 4681
rect 2034 4613 2046 4647
rect 2080 4613 2092 4647
rect 2034 4579 2092 4613
rect 2034 4545 2046 4579
rect 2080 4545 2092 4579
rect 2034 4511 2092 4545
rect 2034 4477 2046 4511
rect 2080 4477 2092 4511
rect 2034 4443 2092 4477
rect 2034 4409 2046 4443
rect 2080 4409 2092 4443
rect 2034 4375 2092 4409
rect 2034 4341 2046 4375
rect 2080 4341 2092 4375
rect 2034 4307 2092 4341
rect 2034 4273 2046 4307
rect 2080 4273 2092 4307
rect 2034 4239 2092 4273
rect 2034 4205 2046 4239
rect 2080 4205 2092 4239
rect 2034 4171 2092 4205
rect 2034 4137 2046 4171
rect 2080 4137 2092 4171
rect 2034 4103 2092 4137
rect 2034 4069 2046 4103
rect 2080 4069 2092 4103
rect 2034 4035 2092 4069
rect 2034 4001 2046 4035
rect 2080 4001 2092 4035
rect 2034 3967 2092 4001
rect 2034 3933 2046 3967
rect 2080 3933 2092 3967
rect 2034 3899 2092 3933
rect 2034 3865 2046 3899
rect 2080 3865 2092 3899
rect 2034 3831 2092 3865
rect 2034 3797 2046 3831
rect 2080 3797 2092 3831
rect 2034 3763 2092 3797
rect 2034 3729 2046 3763
rect 2080 3729 2092 3763
rect 2034 3695 2092 3729
rect 2034 3661 2046 3695
rect 2080 3661 2092 3695
rect 2034 3630 2092 3661
rect 2292 5599 2350 5630
rect 2292 5565 2304 5599
rect 2338 5565 2350 5599
rect 2292 5531 2350 5565
rect 2292 5497 2304 5531
rect 2338 5497 2350 5531
rect 2292 5463 2350 5497
rect 2292 5429 2304 5463
rect 2338 5429 2350 5463
rect 2292 5395 2350 5429
rect 2292 5361 2304 5395
rect 2338 5361 2350 5395
rect 2292 5327 2350 5361
rect 2292 5293 2304 5327
rect 2338 5293 2350 5327
rect 2292 5259 2350 5293
rect 2292 5225 2304 5259
rect 2338 5225 2350 5259
rect 2292 5191 2350 5225
rect 2292 5157 2304 5191
rect 2338 5157 2350 5191
rect 2292 5123 2350 5157
rect 2292 5089 2304 5123
rect 2338 5089 2350 5123
rect 2292 5055 2350 5089
rect 2292 5021 2304 5055
rect 2338 5021 2350 5055
rect 2292 4987 2350 5021
rect 2292 4953 2304 4987
rect 2338 4953 2350 4987
rect 2292 4919 2350 4953
rect 2292 4885 2304 4919
rect 2338 4885 2350 4919
rect 2292 4851 2350 4885
rect 2292 4817 2304 4851
rect 2338 4817 2350 4851
rect 2292 4783 2350 4817
rect 2292 4749 2304 4783
rect 2338 4749 2350 4783
rect 2292 4715 2350 4749
rect 2292 4681 2304 4715
rect 2338 4681 2350 4715
rect 2292 4647 2350 4681
rect 2292 4613 2304 4647
rect 2338 4613 2350 4647
rect 2292 4579 2350 4613
rect 2292 4545 2304 4579
rect 2338 4545 2350 4579
rect 2292 4511 2350 4545
rect 2292 4477 2304 4511
rect 2338 4477 2350 4511
rect 2292 4443 2350 4477
rect 2292 4409 2304 4443
rect 2338 4409 2350 4443
rect 2292 4375 2350 4409
rect 2292 4341 2304 4375
rect 2338 4341 2350 4375
rect 2292 4307 2350 4341
rect 2292 4273 2304 4307
rect 2338 4273 2350 4307
rect 2292 4239 2350 4273
rect 2292 4205 2304 4239
rect 2338 4205 2350 4239
rect 2292 4171 2350 4205
rect 2292 4137 2304 4171
rect 2338 4137 2350 4171
rect 2292 4103 2350 4137
rect 2292 4069 2304 4103
rect 2338 4069 2350 4103
rect 2292 4035 2350 4069
rect 2292 4001 2304 4035
rect 2338 4001 2350 4035
rect 2292 3967 2350 4001
rect 2292 3933 2304 3967
rect 2338 3933 2350 3967
rect 2292 3899 2350 3933
rect 2292 3865 2304 3899
rect 2338 3865 2350 3899
rect 2292 3831 2350 3865
rect 2292 3797 2304 3831
rect 2338 3797 2350 3831
rect 2292 3763 2350 3797
rect 2292 3729 2304 3763
rect 2338 3729 2350 3763
rect 2292 3695 2350 3729
rect 2292 3661 2304 3695
rect 2338 3661 2350 3695
rect 2292 3630 2350 3661
rect 3734 5599 3792 5630
rect 3734 5565 3746 5599
rect 3780 5565 3792 5599
rect 3734 5531 3792 5565
rect 3734 5497 3746 5531
rect 3780 5497 3792 5531
rect 3734 5463 3792 5497
rect 3734 5429 3746 5463
rect 3780 5429 3792 5463
rect 3734 5395 3792 5429
rect 3734 5361 3746 5395
rect 3780 5361 3792 5395
rect 3734 5327 3792 5361
rect 3734 5293 3746 5327
rect 3780 5293 3792 5327
rect 3734 5259 3792 5293
rect 3734 5225 3746 5259
rect 3780 5225 3792 5259
rect 3734 5191 3792 5225
rect 3734 5157 3746 5191
rect 3780 5157 3792 5191
rect 3734 5123 3792 5157
rect 3734 5089 3746 5123
rect 3780 5089 3792 5123
rect 3734 5055 3792 5089
rect 3734 5021 3746 5055
rect 3780 5021 3792 5055
rect 3734 4987 3792 5021
rect 3734 4953 3746 4987
rect 3780 4953 3792 4987
rect 3734 4919 3792 4953
rect 3734 4885 3746 4919
rect 3780 4885 3792 4919
rect 3734 4851 3792 4885
rect 3734 4817 3746 4851
rect 3780 4817 3792 4851
rect 3734 4783 3792 4817
rect 3734 4749 3746 4783
rect 3780 4749 3792 4783
rect 3734 4715 3792 4749
rect 3734 4681 3746 4715
rect 3780 4681 3792 4715
rect 3734 4647 3792 4681
rect 3734 4613 3746 4647
rect 3780 4613 3792 4647
rect 3734 4579 3792 4613
rect 3734 4545 3746 4579
rect 3780 4545 3792 4579
rect 3734 4511 3792 4545
rect 3734 4477 3746 4511
rect 3780 4477 3792 4511
rect 3734 4443 3792 4477
rect 3734 4409 3746 4443
rect 3780 4409 3792 4443
rect 3734 4375 3792 4409
rect 3734 4341 3746 4375
rect 3780 4341 3792 4375
rect 3734 4307 3792 4341
rect 3734 4273 3746 4307
rect 3780 4273 3792 4307
rect 3734 4239 3792 4273
rect 3734 4205 3746 4239
rect 3780 4205 3792 4239
rect 3734 4171 3792 4205
rect 3734 4137 3746 4171
rect 3780 4137 3792 4171
rect 3734 4103 3792 4137
rect 3734 4069 3746 4103
rect 3780 4069 3792 4103
rect 3734 4035 3792 4069
rect 3734 4001 3746 4035
rect 3780 4001 3792 4035
rect 3734 3967 3792 4001
rect 3734 3933 3746 3967
rect 3780 3933 3792 3967
rect 3734 3899 3792 3933
rect 3734 3865 3746 3899
rect 3780 3865 3792 3899
rect 3734 3831 3792 3865
rect 3734 3797 3746 3831
rect 3780 3797 3792 3831
rect 3734 3763 3792 3797
rect 3734 3729 3746 3763
rect 3780 3729 3792 3763
rect 3734 3695 3792 3729
rect 3734 3661 3746 3695
rect 3780 3661 3792 3695
rect 3734 3630 3792 3661
rect 3992 5599 4050 5630
rect 3992 5565 4004 5599
rect 4038 5565 4050 5599
rect 3992 5531 4050 5565
rect 3992 5497 4004 5531
rect 4038 5497 4050 5531
rect 3992 5463 4050 5497
rect 3992 5429 4004 5463
rect 4038 5429 4050 5463
rect 3992 5395 4050 5429
rect 3992 5361 4004 5395
rect 4038 5361 4050 5395
rect 3992 5327 4050 5361
rect 3992 5293 4004 5327
rect 4038 5293 4050 5327
rect 3992 5259 4050 5293
rect 3992 5225 4004 5259
rect 4038 5225 4050 5259
rect 3992 5191 4050 5225
rect 3992 5157 4004 5191
rect 4038 5157 4050 5191
rect 3992 5123 4050 5157
rect 3992 5089 4004 5123
rect 4038 5089 4050 5123
rect 3992 5055 4050 5089
rect 3992 5021 4004 5055
rect 4038 5021 4050 5055
rect 3992 4987 4050 5021
rect 3992 4953 4004 4987
rect 4038 4953 4050 4987
rect 3992 4919 4050 4953
rect 3992 4885 4004 4919
rect 4038 4885 4050 4919
rect 3992 4851 4050 4885
rect 3992 4817 4004 4851
rect 4038 4817 4050 4851
rect 3992 4783 4050 4817
rect 3992 4749 4004 4783
rect 4038 4749 4050 4783
rect 3992 4715 4050 4749
rect 3992 4681 4004 4715
rect 4038 4681 4050 4715
rect 3992 4647 4050 4681
rect 3992 4613 4004 4647
rect 4038 4613 4050 4647
rect 3992 4579 4050 4613
rect 3992 4545 4004 4579
rect 4038 4545 4050 4579
rect 3992 4511 4050 4545
rect 3992 4477 4004 4511
rect 4038 4477 4050 4511
rect 3992 4443 4050 4477
rect 3992 4409 4004 4443
rect 4038 4409 4050 4443
rect 3992 4375 4050 4409
rect 3992 4341 4004 4375
rect 4038 4341 4050 4375
rect 3992 4307 4050 4341
rect 3992 4273 4004 4307
rect 4038 4273 4050 4307
rect 3992 4239 4050 4273
rect 3992 4205 4004 4239
rect 4038 4205 4050 4239
rect 3992 4171 4050 4205
rect 3992 4137 4004 4171
rect 4038 4137 4050 4171
rect 3992 4103 4050 4137
rect 3992 4069 4004 4103
rect 4038 4069 4050 4103
rect 3992 4035 4050 4069
rect 3992 4001 4004 4035
rect 4038 4001 4050 4035
rect 3992 3967 4050 4001
rect 3992 3933 4004 3967
rect 4038 3933 4050 3967
rect 3992 3899 4050 3933
rect 3992 3865 4004 3899
rect 4038 3865 4050 3899
rect 3992 3831 4050 3865
rect 3992 3797 4004 3831
rect 4038 3797 4050 3831
rect 3992 3763 4050 3797
rect 3992 3729 4004 3763
rect 4038 3729 4050 3763
rect 3992 3695 4050 3729
rect 3992 3661 4004 3695
rect 4038 3661 4050 3695
rect 3992 3630 4050 3661
rect 4434 5599 4492 5630
rect 4434 5565 4446 5599
rect 4480 5565 4492 5599
rect 4434 5531 4492 5565
rect 4434 5497 4446 5531
rect 4480 5497 4492 5531
rect 4434 5463 4492 5497
rect 4434 5429 4446 5463
rect 4480 5429 4492 5463
rect 4434 5395 4492 5429
rect 4434 5361 4446 5395
rect 4480 5361 4492 5395
rect 4434 5327 4492 5361
rect 4434 5293 4446 5327
rect 4480 5293 4492 5327
rect 4434 5259 4492 5293
rect 4434 5225 4446 5259
rect 4480 5225 4492 5259
rect 4434 5191 4492 5225
rect 4434 5157 4446 5191
rect 4480 5157 4492 5191
rect 4434 5123 4492 5157
rect 4434 5089 4446 5123
rect 4480 5089 4492 5123
rect 4434 5055 4492 5089
rect 4434 5021 4446 5055
rect 4480 5021 4492 5055
rect 4434 4987 4492 5021
rect 4434 4953 4446 4987
rect 4480 4953 4492 4987
rect 4434 4919 4492 4953
rect 4434 4885 4446 4919
rect 4480 4885 4492 4919
rect 4434 4851 4492 4885
rect 4434 4817 4446 4851
rect 4480 4817 4492 4851
rect 4434 4783 4492 4817
rect 4434 4749 4446 4783
rect 4480 4749 4492 4783
rect 4434 4715 4492 4749
rect 4434 4681 4446 4715
rect 4480 4681 4492 4715
rect 4434 4647 4492 4681
rect 4434 4613 4446 4647
rect 4480 4613 4492 4647
rect 4434 4579 4492 4613
rect 4434 4545 4446 4579
rect 4480 4545 4492 4579
rect 4434 4511 4492 4545
rect 4434 4477 4446 4511
rect 4480 4477 4492 4511
rect 4434 4443 4492 4477
rect 4434 4409 4446 4443
rect 4480 4409 4492 4443
rect 4434 4375 4492 4409
rect 4434 4341 4446 4375
rect 4480 4341 4492 4375
rect 4434 4307 4492 4341
rect 4434 4273 4446 4307
rect 4480 4273 4492 4307
rect 4434 4239 4492 4273
rect 4434 4205 4446 4239
rect 4480 4205 4492 4239
rect 4434 4171 4492 4205
rect 4434 4137 4446 4171
rect 4480 4137 4492 4171
rect 4434 4103 4492 4137
rect 4434 4069 4446 4103
rect 4480 4069 4492 4103
rect 4434 4035 4492 4069
rect 4434 4001 4446 4035
rect 4480 4001 4492 4035
rect 4434 3967 4492 4001
rect 4434 3933 4446 3967
rect 4480 3933 4492 3967
rect 4434 3899 4492 3933
rect 4434 3865 4446 3899
rect 4480 3865 4492 3899
rect 4434 3831 4492 3865
rect 4434 3797 4446 3831
rect 4480 3797 4492 3831
rect 4434 3763 4492 3797
rect 4434 3729 4446 3763
rect 4480 3729 4492 3763
rect 4434 3695 4492 3729
rect 4434 3661 4446 3695
rect 4480 3661 4492 3695
rect 4434 3630 4492 3661
rect 4692 5599 4750 5630
rect 4692 5565 4704 5599
rect 4738 5565 4750 5599
rect 4692 5531 4750 5565
rect 4692 5497 4704 5531
rect 4738 5497 4750 5531
rect 4692 5463 4750 5497
rect 4692 5429 4704 5463
rect 4738 5429 4750 5463
rect 4692 5395 4750 5429
rect 4692 5361 4704 5395
rect 4738 5361 4750 5395
rect 4692 5327 4750 5361
rect 4692 5293 4704 5327
rect 4738 5293 4750 5327
rect 4692 5259 4750 5293
rect 4692 5225 4704 5259
rect 4738 5225 4750 5259
rect 4692 5191 4750 5225
rect 4692 5157 4704 5191
rect 4738 5157 4750 5191
rect 4692 5123 4750 5157
rect 4692 5089 4704 5123
rect 4738 5089 4750 5123
rect 4692 5055 4750 5089
rect 4692 5021 4704 5055
rect 4738 5021 4750 5055
rect 4692 4987 4750 5021
rect 4692 4953 4704 4987
rect 4738 4953 4750 4987
rect 4692 4919 4750 4953
rect 4692 4885 4704 4919
rect 4738 4885 4750 4919
rect 4692 4851 4750 4885
rect 4692 4817 4704 4851
rect 4738 4817 4750 4851
rect 4692 4783 4750 4817
rect 4692 4749 4704 4783
rect 4738 4749 4750 4783
rect 4692 4715 4750 4749
rect 4692 4681 4704 4715
rect 4738 4681 4750 4715
rect 4692 4647 4750 4681
rect 4692 4613 4704 4647
rect 4738 4613 4750 4647
rect 4692 4579 4750 4613
rect 4692 4545 4704 4579
rect 4738 4545 4750 4579
rect 4692 4511 4750 4545
rect 4692 4477 4704 4511
rect 4738 4477 4750 4511
rect 4692 4443 4750 4477
rect 4692 4409 4704 4443
rect 4738 4409 4750 4443
rect 4692 4375 4750 4409
rect 4692 4341 4704 4375
rect 4738 4341 4750 4375
rect 4692 4307 4750 4341
rect 4692 4273 4704 4307
rect 4738 4273 4750 4307
rect 4692 4239 4750 4273
rect 4692 4205 4704 4239
rect 4738 4205 4750 4239
rect 4692 4171 4750 4205
rect 4692 4137 4704 4171
rect 4738 4137 4750 4171
rect 4692 4103 4750 4137
rect 4692 4069 4704 4103
rect 4738 4069 4750 4103
rect 4692 4035 4750 4069
rect 4692 4001 4704 4035
rect 4738 4001 4750 4035
rect 4692 3967 4750 4001
rect 4692 3933 4704 3967
rect 4738 3933 4750 3967
rect 4692 3899 4750 3933
rect 4692 3865 4704 3899
rect 4738 3865 4750 3899
rect 4692 3831 4750 3865
rect 4692 3797 4704 3831
rect 4738 3797 4750 3831
rect 4692 3763 4750 3797
rect 4692 3729 4704 3763
rect 4738 3729 4750 3763
rect 4692 3695 4750 3729
rect 4692 3661 4704 3695
rect 4738 3661 4750 3695
rect 4692 3630 4750 3661
rect 5134 5599 5192 5630
rect 5134 5565 5146 5599
rect 5180 5565 5192 5599
rect 5134 5531 5192 5565
rect 5134 5497 5146 5531
rect 5180 5497 5192 5531
rect 5134 5463 5192 5497
rect 5134 5429 5146 5463
rect 5180 5429 5192 5463
rect 5134 5395 5192 5429
rect 5134 5361 5146 5395
rect 5180 5361 5192 5395
rect 5134 5327 5192 5361
rect 5134 5293 5146 5327
rect 5180 5293 5192 5327
rect 5134 5259 5192 5293
rect 5134 5225 5146 5259
rect 5180 5225 5192 5259
rect 5134 5191 5192 5225
rect 5134 5157 5146 5191
rect 5180 5157 5192 5191
rect 5134 5123 5192 5157
rect 5134 5089 5146 5123
rect 5180 5089 5192 5123
rect 5134 5055 5192 5089
rect 5134 5021 5146 5055
rect 5180 5021 5192 5055
rect 5134 4987 5192 5021
rect 5134 4953 5146 4987
rect 5180 4953 5192 4987
rect 5134 4919 5192 4953
rect 5134 4885 5146 4919
rect 5180 4885 5192 4919
rect 5134 4851 5192 4885
rect 5134 4817 5146 4851
rect 5180 4817 5192 4851
rect 5134 4783 5192 4817
rect 5134 4749 5146 4783
rect 5180 4749 5192 4783
rect 5134 4715 5192 4749
rect 5134 4681 5146 4715
rect 5180 4681 5192 4715
rect 5134 4647 5192 4681
rect 5134 4613 5146 4647
rect 5180 4613 5192 4647
rect 5134 4579 5192 4613
rect 5134 4545 5146 4579
rect 5180 4545 5192 4579
rect 5134 4511 5192 4545
rect 5134 4477 5146 4511
rect 5180 4477 5192 4511
rect 5134 4443 5192 4477
rect 5134 4409 5146 4443
rect 5180 4409 5192 4443
rect 5134 4375 5192 4409
rect 5134 4341 5146 4375
rect 5180 4341 5192 4375
rect 5134 4307 5192 4341
rect 5134 4273 5146 4307
rect 5180 4273 5192 4307
rect 5134 4239 5192 4273
rect 5134 4205 5146 4239
rect 5180 4205 5192 4239
rect 5134 4171 5192 4205
rect 5134 4137 5146 4171
rect 5180 4137 5192 4171
rect 5134 4103 5192 4137
rect 5134 4069 5146 4103
rect 5180 4069 5192 4103
rect 5134 4035 5192 4069
rect 5134 4001 5146 4035
rect 5180 4001 5192 4035
rect 5134 3967 5192 4001
rect 5134 3933 5146 3967
rect 5180 3933 5192 3967
rect 5134 3899 5192 3933
rect 5134 3865 5146 3899
rect 5180 3865 5192 3899
rect 5134 3831 5192 3865
rect 5134 3797 5146 3831
rect 5180 3797 5192 3831
rect 5134 3763 5192 3797
rect 5134 3729 5146 3763
rect 5180 3729 5192 3763
rect 5134 3695 5192 3729
rect 5134 3661 5146 3695
rect 5180 3661 5192 3695
rect 5134 3630 5192 3661
rect 5392 5599 5450 5630
rect 5392 5565 5404 5599
rect 5438 5565 5450 5599
rect 5392 5531 5450 5565
rect 5392 5497 5404 5531
rect 5438 5497 5450 5531
rect 5392 5463 5450 5497
rect 5392 5429 5404 5463
rect 5438 5429 5450 5463
rect 5392 5395 5450 5429
rect 5392 5361 5404 5395
rect 5438 5361 5450 5395
rect 5392 5327 5450 5361
rect 5392 5293 5404 5327
rect 5438 5293 5450 5327
rect 5392 5259 5450 5293
rect 5392 5225 5404 5259
rect 5438 5225 5450 5259
rect 5392 5191 5450 5225
rect 5392 5157 5404 5191
rect 5438 5157 5450 5191
rect 5392 5123 5450 5157
rect 5392 5089 5404 5123
rect 5438 5089 5450 5123
rect 5392 5055 5450 5089
rect 5392 5021 5404 5055
rect 5438 5021 5450 5055
rect 5392 4987 5450 5021
rect 5392 4953 5404 4987
rect 5438 4953 5450 4987
rect 5392 4919 5450 4953
rect 5392 4885 5404 4919
rect 5438 4885 5450 4919
rect 5392 4851 5450 4885
rect 5392 4817 5404 4851
rect 5438 4817 5450 4851
rect 5392 4783 5450 4817
rect 5392 4749 5404 4783
rect 5438 4749 5450 4783
rect 5392 4715 5450 4749
rect 5392 4681 5404 4715
rect 5438 4681 5450 4715
rect 5392 4647 5450 4681
rect 5392 4613 5404 4647
rect 5438 4613 5450 4647
rect 5392 4579 5450 4613
rect 5392 4545 5404 4579
rect 5438 4545 5450 4579
rect 5392 4511 5450 4545
rect 5392 4477 5404 4511
rect 5438 4477 5450 4511
rect 5392 4443 5450 4477
rect 5392 4409 5404 4443
rect 5438 4409 5450 4443
rect 5392 4375 5450 4409
rect 5392 4341 5404 4375
rect 5438 4341 5450 4375
rect 5392 4307 5450 4341
rect 5392 4273 5404 4307
rect 5438 4273 5450 4307
rect 5392 4239 5450 4273
rect 5392 4205 5404 4239
rect 5438 4205 5450 4239
rect 5392 4171 5450 4205
rect 5392 4137 5404 4171
rect 5438 4137 5450 4171
rect 5392 4103 5450 4137
rect 5392 4069 5404 4103
rect 5438 4069 5450 4103
rect 5392 4035 5450 4069
rect 5392 4001 5404 4035
rect 5438 4001 5450 4035
rect 5392 3967 5450 4001
rect 5392 3933 5404 3967
rect 5438 3933 5450 3967
rect 5392 3899 5450 3933
rect 5392 3865 5404 3899
rect 5438 3865 5450 3899
rect 5392 3831 5450 3865
rect 5392 3797 5404 3831
rect 5438 3797 5450 3831
rect 5392 3763 5450 3797
rect 5392 3729 5404 3763
rect 5438 3729 5450 3763
rect 5392 3695 5450 3729
rect 5392 3661 5404 3695
rect 5438 3661 5450 3695
rect 5392 3630 5450 3661
rect 5834 5599 5892 5630
rect 5834 5565 5846 5599
rect 5880 5565 5892 5599
rect 5834 5531 5892 5565
rect 5834 5497 5846 5531
rect 5880 5497 5892 5531
rect 5834 5463 5892 5497
rect 5834 5429 5846 5463
rect 5880 5429 5892 5463
rect 5834 5395 5892 5429
rect 5834 5361 5846 5395
rect 5880 5361 5892 5395
rect 5834 5327 5892 5361
rect 5834 5293 5846 5327
rect 5880 5293 5892 5327
rect 5834 5259 5892 5293
rect 5834 5225 5846 5259
rect 5880 5225 5892 5259
rect 5834 5191 5892 5225
rect 5834 5157 5846 5191
rect 5880 5157 5892 5191
rect 5834 5123 5892 5157
rect 5834 5089 5846 5123
rect 5880 5089 5892 5123
rect 5834 5055 5892 5089
rect 5834 5021 5846 5055
rect 5880 5021 5892 5055
rect 5834 4987 5892 5021
rect 5834 4953 5846 4987
rect 5880 4953 5892 4987
rect 5834 4919 5892 4953
rect 5834 4885 5846 4919
rect 5880 4885 5892 4919
rect 5834 4851 5892 4885
rect 5834 4817 5846 4851
rect 5880 4817 5892 4851
rect 5834 4783 5892 4817
rect 5834 4749 5846 4783
rect 5880 4749 5892 4783
rect 5834 4715 5892 4749
rect 5834 4681 5846 4715
rect 5880 4681 5892 4715
rect 5834 4647 5892 4681
rect 5834 4613 5846 4647
rect 5880 4613 5892 4647
rect 5834 4579 5892 4613
rect 5834 4545 5846 4579
rect 5880 4545 5892 4579
rect 5834 4511 5892 4545
rect 5834 4477 5846 4511
rect 5880 4477 5892 4511
rect 5834 4443 5892 4477
rect 5834 4409 5846 4443
rect 5880 4409 5892 4443
rect 5834 4375 5892 4409
rect 5834 4341 5846 4375
rect 5880 4341 5892 4375
rect 5834 4307 5892 4341
rect 5834 4273 5846 4307
rect 5880 4273 5892 4307
rect 5834 4239 5892 4273
rect 5834 4205 5846 4239
rect 5880 4205 5892 4239
rect 5834 4171 5892 4205
rect 5834 4137 5846 4171
rect 5880 4137 5892 4171
rect 5834 4103 5892 4137
rect 5834 4069 5846 4103
rect 5880 4069 5892 4103
rect 5834 4035 5892 4069
rect 5834 4001 5846 4035
rect 5880 4001 5892 4035
rect 5834 3967 5892 4001
rect 5834 3933 5846 3967
rect 5880 3933 5892 3967
rect 5834 3899 5892 3933
rect 5834 3865 5846 3899
rect 5880 3865 5892 3899
rect 5834 3831 5892 3865
rect 5834 3797 5846 3831
rect 5880 3797 5892 3831
rect 5834 3763 5892 3797
rect 5834 3729 5846 3763
rect 5880 3729 5892 3763
rect 5834 3695 5892 3729
rect 5834 3661 5846 3695
rect 5880 3661 5892 3695
rect 5834 3630 5892 3661
rect 6092 5599 6150 5630
rect 6092 5565 6104 5599
rect 6138 5565 6150 5599
rect 6092 5531 6150 5565
rect 6092 5497 6104 5531
rect 6138 5497 6150 5531
rect 6092 5463 6150 5497
rect 6092 5429 6104 5463
rect 6138 5429 6150 5463
rect 6092 5395 6150 5429
rect 6092 5361 6104 5395
rect 6138 5361 6150 5395
rect 6092 5327 6150 5361
rect 6092 5293 6104 5327
rect 6138 5293 6150 5327
rect 6092 5259 6150 5293
rect 6092 5225 6104 5259
rect 6138 5225 6150 5259
rect 6092 5191 6150 5225
rect 6092 5157 6104 5191
rect 6138 5157 6150 5191
rect 6092 5123 6150 5157
rect 6092 5089 6104 5123
rect 6138 5089 6150 5123
rect 6092 5055 6150 5089
rect 6092 5021 6104 5055
rect 6138 5021 6150 5055
rect 6092 4987 6150 5021
rect 6092 4953 6104 4987
rect 6138 4953 6150 4987
rect 6092 4919 6150 4953
rect 6092 4885 6104 4919
rect 6138 4885 6150 4919
rect 6092 4851 6150 4885
rect 6092 4817 6104 4851
rect 6138 4817 6150 4851
rect 6092 4783 6150 4817
rect 6092 4749 6104 4783
rect 6138 4749 6150 4783
rect 6092 4715 6150 4749
rect 6092 4681 6104 4715
rect 6138 4681 6150 4715
rect 6092 4647 6150 4681
rect 6092 4613 6104 4647
rect 6138 4613 6150 4647
rect 6092 4579 6150 4613
rect 6092 4545 6104 4579
rect 6138 4545 6150 4579
rect 6092 4511 6150 4545
rect 6092 4477 6104 4511
rect 6138 4477 6150 4511
rect 6092 4443 6150 4477
rect 6092 4409 6104 4443
rect 6138 4409 6150 4443
rect 6092 4375 6150 4409
rect 6092 4341 6104 4375
rect 6138 4341 6150 4375
rect 6092 4307 6150 4341
rect 6092 4273 6104 4307
rect 6138 4273 6150 4307
rect 6092 4239 6150 4273
rect 6092 4205 6104 4239
rect 6138 4205 6150 4239
rect 6092 4171 6150 4205
rect 6092 4137 6104 4171
rect 6138 4137 6150 4171
rect 6092 4103 6150 4137
rect 6092 4069 6104 4103
rect 6138 4069 6150 4103
rect 6092 4035 6150 4069
rect 6092 4001 6104 4035
rect 6138 4001 6150 4035
rect 6092 3967 6150 4001
rect 6092 3933 6104 3967
rect 6138 3933 6150 3967
rect 6092 3899 6150 3933
rect 6092 3865 6104 3899
rect 6138 3865 6150 3899
rect 6092 3831 6150 3865
rect 6092 3797 6104 3831
rect 6138 3797 6150 3831
rect 6092 3763 6150 3797
rect 6092 3729 6104 3763
rect 6138 3729 6150 3763
rect 6092 3695 6150 3729
rect 6092 3661 6104 3695
rect 6138 3661 6150 3695
rect 6092 3630 6150 3661
rect 6534 5599 6592 5630
rect 6534 5565 6546 5599
rect 6580 5565 6592 5599
rect 6534 5531 6592 5565
rect 6534 5497 6546 5531
rect 6580 5497 6592 5531
rect 6534 5463 6592 5497
rect 6534 5429 6546 5463
rect 6580 5429 6592 5463
rect 6534 5395 6592 5429
rect 6534 5361 6546 5395
rect 6580 5361 6592 5395
rect 6534 5327 6592 5361
rect 6534 5293 6546 5327
rect 6580 5293 6592 5327
rect 6534 5259 6592 5293
rect 6534 5225 6546 5259
rect 6580 5225 6592 5259
rect 6534 5191 6592 5225
rect 6534 5157 6546 5191
rect 6580 5157 6592 5191
rect 6534 5123 6592 5157
rect 6534 5089 6546 5123
rect 6580 5089 6592 5123
rect 6534 5055 6592 5089
rect 6534 5021 6546 5055
rect 6580 5021 6592 5055
rect 6534 4987 6592 5021
rect 6534 4953 6546 4987
rect 6580 4953 6592 4987
rect 6534 4919 6592 4953
rect 6534 4885 6546 4919
rect 6580 4885 6592 4919
rect 6534 4851 6592 4885
rect 6534 4817 6546 4851
rect 6580 4817 6592 4851
rect 6534 4783 6592 4817
rect 6534 4749 6546 4783
rect 6580 4749 6592 4783
rect 6534 4715 6592 4749
rect 6534 4681 6546 4715
rect 6580 4681 6592 4715
rect 6534 4647 6592 4681
rect 6534 4613 6546 4647
rect 6580 4613 6592 4647
rect 6534 4579 6592 4613
rect 6534 4545 6546 4579
rect 6580 4545 6592 4579
rect 6534 4511 6592 4545
rect 6534 4477 6546 4511
rect 6580 4477 6592 4511
rect 6534 4443 6592 4477
rect 6534 4409 6546 4443
rect 6580 4409 6592 4443
rect 6534 4375 6592 4409
rect 6534 4341 6546 4375
rect 6580 4341 6592 4375
rect 6534 4307 6592 4341
rect 6534 4273 6546 4307
rect 6580 4273 6592 4307
rect 6534 4239 6592 4273
rect 6534 4205 6546 4239
rect 6580 4205 6592 4239
rect 6534 4171 6592 4205
rect 6534 4137 6546 4171
rect 6580 4137 6592 4171
rect 6534 4103 6592 4137
rect 6534 4069 6546 4103
rect 6580 4069 6592 4103
rect 6534 4035 6592 4069
rect 6534 4001 6546 4035
rect 6580 4001 6592 4035
rect 6534 3967 6592 4001
rect 6534 3933 6546 3967
rect 6580 3933 6592 3967
rect 6534 3899 6592 3933
rect 6534 3865 6546 3899
rect 6580 3865 6592 3899
rect 6534 3831 6592 3865
rect 6534 3797 6546 3831
rect 6580 3797 6592 3831
rect 6534 3763 6592 3797
rect 6534 3729 6546 3763
rect 6580 3729 6592 3763
rect 6534 3695 6592 3729
rect 6534 3661 6546 3695
rect 6580 3661 6592 3695
rect 6534 3630 6592 3661
rect 6792 5599 6850 5630
rect 6792 5565 6804 5599
rect 6838 5565 6850 5599
rect 6792 5531 6850 5565
rect 6792 5497 6804 5531
rect 6838 5497 6850 5531
rect 6792 5463 6850 5497
rect 6792 5429 6804 5463
rect 6838 5429 6850 5463
rect 6792 5395 6850 5429
rect 6792 5361 6804 5395
rect 6838 5361 6850 5395
rect 6792 5327 6850 5361
rect 6792 5293 6804 5327
rect 6838 5293 6850 5327
rect 6792 5259 6850 5293
rect 6792 5225 6804 5259
rect 6838 5225 6850 5259
rect 6792 5191 6850 5225
rect 6792 5157 6804 5191
rect 6838 5157 6850 5191
rect 6792 5123 6850 5157
rect 6792 5089 6804 5123
rect 6838 5089 6850 5123
rect 6792 5055 6850 5089
rect 6792 5021 6804 5055
rect 6838 5021 6850 5055
rect 6792 4987 6850 5021
rect 6792 4953 6804 4987
rect 6838 4953 6850 4987
rect 6792 4919 6850 4953
rect 6792 4885 6804 4919
rect 6838 4885 6850 4919
rect 6792 4851 6850 4885
rect 6792 4817 6804 4851
rect 6838 4817 6850 4851
rect 6792 4783 6850 4817
rect 6792 4749 6804 4783
rect 6838 4749 6850 4783
rect 6792 4715 6850 4749
rect 6792 4681 6804 4715
rect 6838 4681 6850 4715
rect 6792 4647 6850 4681
rect 6792 4613 6804 4647
rect 6838 4613 6850 4647
rect 6792 4579 6850 4613
rect 6792 4545 6804 4579
rect 6838 4545 6850 4579
rect 6792 4511 6850 4545
rect 6792 4477 6804 4511
rect 6838 4477 6850 4511
rect 6792 4443 6850 4477
rect 6792 4409 6804 4443
rect 6838 4409 6850 4443
rect 6792 4375 6850 4409
rect 6792 4341 6804 4375
rect 6838 4341 6850 4375
rect 6792 4307 6850 4341
rect 6792 4273 6804 4307
rect 6838 4273 6850 4307
rect 6792 4239 6850 4273
rect 6792 4205 6804 4239
rect 6838 4205 6850 4239
rect 6792 4171 6850 4205
rect 6792 4137 6804 4171
rect 6838 4137 6850 4171
rect 6792 4103 6850 4137
rect 6792 4069 6804 4103
rect 6838 4069 6850 4103
rect 6792 4035 6850 4069
rect 6792 4001 6804 4035
rect 6838 4001 6850 4035
rect 6792 3967 6850 4001
rect 6792 3933 6804 3967
rect 6838 3933 6850 3967
rect 6792 3899 6850 3933
rect 6792 3865 6804 3899
rect 6838 3865 6850 3899
rect 6792 3831 6850 3865
rect 6792 3797 6804 3831
rect 6838 3797 6850 3831
rect 6792 3763 6850 3797
rect 6792 3729 6804 3763
rect 6838 3729 6850 3763
rect 6792 3695 6850 3729
rect 6792 3661 6804 3695
rect 6838 3661 6850 3695
rect 6792 3630 6850 3661
rect 7234 5599 7292 5630
rect 7234 5565 7246 5599
rect 7280 5565 7292 5599
rect 7234 5531 7292 5565
rect 7234 5497 7246 5531
rect 7280 5497 7292 5531
rect 7234 5463 7292 5497
rect 7234 5429 7246 5463
rect 7280 5429 7292 5463
rect 7234 5395 7292 5429
rect 7234 5361 7246 5395
rect 7280 5361 7292 5395
rect 7234 5327 7292 5361
rect 7234 5293 7246 5327
rect 7280 5293 7292 5327
rect 7234 5259 7292 5293
rect 7234 5225 7246 5259
rect 7280 5225 7292 5259
rect 7234 5191 7292 5225
rect 7234 5157 7246 5191
rect 7280 5157 7292 5191
rect 7234 5123 7292 5157
rect 7234 5089 7246 5123
rect 7280 5089 7292 5123
rect 7234 5055 7292 5089
rect 7234 5021 7246 5055
rect 7280 5021 7292 5055
rect 7234 4987 7292 5021
rect 7234 4953 7246 4987
rect 7280 4953 7292 4987
rect 7234 4919 7292 4953
rect 7234 4885 7246 4919
rect 7280 4885 7292 4919
rect 7234 4851 7292 4885
rect 7234 4817 7246 4851
rect 7280 4817 7292 4851
rect 7234 4783 7292 4817
rect 7234 4749 7246 4783
rect 7280 4749 7292 4783
rect 7234 4715 7292 4749
rect 7234 4681 7246 4715
rect 7280 4681 7292 4715
rect 7234 4647 7292 4681
rect 7234 4613 7246 4647
rect 7280 4613 7292 4647
rect 7234 4579 7292 4613
rect 7234 4545 7246 4579
rect 7280 4545 7292 4579
rect 7234 4511 7292 4545
rect 7234 4477 7246 4511
rect 7280 4477 7292 4511
rect 7234 4443 7292 4477
rect 7234 4409 7246 4443
rect 7280 4409 7292 4443
rect 7234 4375 7292 4409
rect 7234 4341 7246 4375
rect 7280 4341 7292 4375
rect 7234 4307 7292 4341
rect 7234 4273 7246 4307
rect 7280 4273 7292 4307
rect 7234 4239 7292 4273
rect 7234 4205 7246 4239
rect 7280 4205 7292 4239
rect 7234 4171 7292 4205
rect 7234 4137 7246 4171
rect 7280 4137 7292 4171
rect 7234 4103 7292 4137
rect 7234 4069 7246 4103
rect 7280 4069 7292 4103
rect 7234 4035 7292 4069
rect 7234 4001 7246 4035
rect 7280 4001 7292 4035
rect 7234 3967 7292 4001
rect 7234 3933 7246 3967
rect 7280 3933 7292 3967
rect 7234 3899 7292 3933
rect 7234 3865 7246 3899
rect 7280 3865 7292 3899
rect 7234 3831 7292 3865
rect 7234 3797 7246 3831
rect 7280 3797 7292 3831
rect 7234 3763 7292 3797
rect 7234 3729 7246 3763
rect 7280 3729 7292 3763
rect 7234 3695 7292 3729
rect 7234 3661 7246 3695
rect 7280 3661 7292 3695
rect 7234 3630 7292 3661
rect 7492 5599 7550 5630
rect 7492 5565 7504 5599
rect 7538 5565 7550 5599
rect 7492 5531 7550 5565
rect 7492 5497 7504 5531
rect 7538 5497 7550 5531
rect 7492 5463 7550 5497
rect 7492 5429 7504 5463
rect 7538 5429 7550 5463
rect 7492 5395 7550 5429
rect 7492 5361 7504 5395
rect 7538 5361 7550 5395
rect 7492 5327 7550 5361
rect 7492 5293 7504 5327
rect 7538 5293 7550 5327
rect 7492 5259 7550 5293
rect 7492 5225 7504 5259
rect 7538 5225 7550 5259
rect 7492 5191 7550 5225
rect 7492 5157 7504 5191
rect 7538 5157 7550 5191
rect 7492 5123 7550 5157
rect 7492 5089 7504 5123
rect 7538 5089 7550 5123
rect 7492 5055 7550 5089
rect 7492 5021 7504 5055
rect 7538 5021 7550 5055
rect 7492 4987 7550 5021
rect 7492 4953 7504 4987
rect 7538 4953 7550 4987
rect 7492 4919 7550 4953
rect 7492 4885 7504 4919
rect 7538 4885 7550 4919
rect 7492 4851 7550 4885
rect 7492 4817 7504 4851
rect 7538 4817 7550 4851
rect 7492 4783 7550 4817
rect 7492 4749 7504 4783
rect 7538 4749 7550 4783
rect 7492 4715 7550 4749
rect 7492 4681 7504 4715
rect 7538 4681 7550 4715
rect 7492 4647 7550 4681
rect 7492 4613 7504 4647
rect 7538 4613 7550 4647
rect 7492 4579 7550 4613
rect 7492 4545 7504 4579
rect 7538 4545 7550 4579
rect 7492 4511 7550 4545
rect 7492 4477 7504 4511
rect 7538 4477 7550 4511
rect 7492 4443 7550 4477
rect 7492 4409 7504 4443
rect 7538 4409 7550 4443
rect 7492 4375 7550 4409
rect 7492 4341 7504 4375
rect 7538 4341 7550 4375
rect 7492 4307 7550 4341
rect 7492 4273 7504 4307
rect 7538 4273 7550 4307
rect 7492 4239 7550 4273
rect 7492 4205 7504 4239
rect 7538 4205 7550 4239
rect 7492 4171 7550 4205
rect 7492 4137 7504 4171
rect 7538 4137 7550 4171
rect 7492 4103 7550 4137
rect 7492 4069 7504 4103
rect 7538 4069 7550 4103
rect 7492 4035 7550 4069
rect 7492 4001 7504 4035
rect 7538 4001 7550 4035
rect 7492 3967 7550 4001
rect 7492 3933 7504 3967
rect 7538 3933 7550 3967
rect 7492 3899 7550 3933
rect 7492 3865 7504 3899
rect 7538 3865 7550 3899
rect 7492 3831 7550 3865
rect 7492 3797 7504 3831
rect 7538 3797 7550 3831
rect 7492 3763 7550 3797
rect 7492 3729 7504 3763
rect 7538 3729 7550 3763
rect 7492 3695 7550 3729
rect 7492 3661 7504 3695
rect 7538 3661 7550 3695
rect 7492 3630 7550 3661
rect 7934 5599 7992 5630
rect 7934 5565 7946 5599
rect 7980 5565 7992 5599
rect 7934 5531 7992 5565
rect 7934 5497 7946 5531
rect 7980 5497 7992 5531
rect 7934 5463 7992 5497
rect 7934 5429 7946 5463
rect 7980 5429 7992 5463
rect 7934 5395 7992 5429
rect 7934 5361 7946 5395
rect 7980 5361 7992 5395
rect 7934 5327 7992 5361
rect 7934 5293 7946 5327
rect 7980 5293 7992 5327
rect 7934 5259 7992 5293
rect 7934 5225 7946 5259
rect 7980 5225 7992 5259
rect 7934 5191 7992 5225
rect 7934 5157 7946 5191
rect 7980 5157 7992 5191
rect 7934 5123 7992 5157
rect 7934 5089 7946 5123
rect 7980 5089 7992 5123
rect 7934 5055 7992 5089
rect 7934 5021 7946 5055
rect 7980 5021 7992 5055
rect 7934 4987 7992 5021
rect 7934 4953 7946 4987
rect 7980 4953 7992 4987
rect 7934 4919 7992 4953
rect 7934 4885 7946 4919
rect 7980 4885 7992 4919
rect 7934 4851 7992 4885
rect 7934 4817 7946 4851
rect 7980 4817 7992 4851
rect 7934 4783 7992 4817
rect 7934 4749 7946 4783
rect 7980 4749 7992 4783
rect 7934 4715 7992 4749
rect 7934 4681 7946 4715
rect 7980 4681 7992 4715
rect 7934 4647 7992 4681
rect 7934 4613 7946 4647
rect 7980 4613 7992 4647
rect 7934 4579 7992 4613
rect 7934 4545 7946 4579
rect 7980 4545 7992 4579
rect 7934 4511 7992 4545
rect 7934 4477 7946 4511
rect 7980 4477 7992 4511
rect 7934 4443 7992 4477
rect 7934 4409 7946 4443
rect 7980 4409 7992 4443
rect 7934 4375 7992 4409
rect 7934 4341 7946 4375
rect 7980 4341 7992 4375
rect 7934 4307 7992 4341
rect 7934 4273 7946 4307
rect 7980 4273 7992 4307
rect 7934 4239 7992 4273
rect 7934 4205 7946 4239
rect 7980 4205 7992 4239
rect 7934 4171 7992 4205
rect 7934 4137 7946 4171
rect 7980 4137 7992 4171
rect 7934 4103 7992 4137
rect 7934 4069 7946 4103
rect 7980 4069 7992 4103
rect 7934 4035 7992 4069
rect 7934 4001 7946 4035
rect 7980 4001 7992 4035
rect 7934 3967 7992 4001
rect 7934 3933 7946 3967
rect 7980 3933 7992 3967
rect 7934 3899 7992 3933
rect 7934 3865 7946 3899
rect 7980 3865 7992 3899
rect 7934 3831 7992 3865
rect 7934 3797 7946 3831
rect 7980 3797 7992 3831
rect 7934 3763 7992 3797
rect 7934 3729 7946 3763
rect 7980 3729 7992 3763
rect 7934 3695 7992 3729
rect 7934 3661 7946 3695
rect 7980 3661 7992 3695
rect 7934 3630 7992 3661
rect 8192 5599 8250 5630
rect 8192 5565 8204 5599
rect 8238 5565 8250 5599
rect 8192 5531 8250 5565
rect 8192 5497 8204 5531
rect 8238 5497 8250 5531
rect 8192 5463 8250 5497
rect 8192 5429 8204 5463
rect 8238 5429 8250 5463
rect 8192 5395 8250 5429
rect 8192 5361 8204 5395
rect 8238 5361 8250 5395
rect 8192 5327 8250 5361
rect 8192 5293 8204 5327
rect 8238 5293 8250 5327
rect 8192 5259 8250 5293
rect 8192 5225 8204 5259
rect 8238 5225 8250 5259
rect 8192 5191 8250 5225
rect 8192 5157 8204 5191
rect 8238 5157 8250 5191
rect 8192 5123 8250 5157
rect 8192 5089 8204 5123
rect 8238 5089 8250 5123
rect 8192 5055 8250 5089
rect 8192 5021 8204 5055
rect 8238 5021 8250 5055
rect 8192 4987 8250 5021
rect 8192 4953 8204 4987
rect 8238 4953 8250 4987
rect 8192 4919 8250 4953
rect 8192 4885 8204 4919
rect 8238 4885 8250 4919
rect 8192 4851 8250 4885
rect 8192 4817 8204 4851
rect 8238 4817 8250 4851
rect 8192 4783 8250 4817
rect 8192 4749 8204 4783
rect 8238 4749 8250 4783
rect 8192 4715 8250 4749
rect 8192 4681 8204 4715
rect 8238 4681 8250 4715
rect 8192 4647 8250 4681
rect 8192 4613 8204 4647
rect 8238 4613 8250 4647
rect 8192 4579 8250 4613
rect 8192 4545 8204 4579
rect 8238 4545 8250 4579
rect 8192 4511 8250 4545
rect 8192 4477 8204 4511
rect 8238 4477 8250 4511
rect 8192 4443 8250 4477
rect 8192 4409 8204 4443
rect 8238 4409 8250 4443
rect 8192 4375 8250 4409
rect 8192 4341 8204 4375
rect 8238 4341 8250 4375
rect 8192 4307 8250 4341
rect 8192 4273 8204 4307
rect 8238 4273 8250 4307
rect 8192 4239 8250 4273
rect 8192 4205 8204 4239
rect 8238 4205 8250 4239
rect 8192 4171 8250 4205
rect 8192 4137 8204 4171
rect 8238 4137 8250 4171
rect 8192 4103 8250 4137
rect 8192 4069 8204 4103
rect 8238 4069 8250 4103
rect 8192 4035 8250 4069
rect 8192 4001 8204 4035
rect 8238 4001 8250 4035
rect 8192 3967 8250 4001
rect 8192 3933 8204 3967
rect 8238 3933 8250 3967
rect 8192 3899 8250 3933
rect 8192 3865 8204 3899
rect 8238 3865 8250 3899
rect 8192 3831 8250 3865
rect 8192 3797 8204 3831
rect 8238 3797 8250 3831
rect 8192 3763 8250 3797
rect 8192 3729 8204 3763
rect 8238 3729 8250 3763
rect 8192 3695 8250 3729
rect 8192 3661 8204 3695
rect 8238 3661 8250 3695
rect 8192 3630 8250 3661
rect 8634 5599 8692 5630
rect 8634 5565 8646 5599
rect 8680 5565 8692 5599
rect 8634 5531 8692 5565
rect 8634 5497 8646 5531
rect 8680 5497 8692 5531
rect 8634 5463 8692 5497
rect 8634 5429 8646 5463
rect 8680 5429 8692 5463
rect 8634 5395 8692 5429
rect 8634 5361 8646 5395
rect 8680 5361 8692 5395
rect 8634 5327 8692 5361
rect 8634 5293 8646 5327
rect 8680 5293 8692 5327
rect 8634 5259 8692 5293
rect 8634 5225 8646 5259
rect 8680 5225 8692 5259
rect 8634 5191 8692 5225
rect 8634 5157 8646 5191
rect 8680 5157 8692 5191
rect 8634 5123 8692 5157
rect 8634 5089 8646 5123
rect 8680 5089 8692 5123
rect 8634 5055 8692 5089
rect 8634 5021 8646 5055
rect 8680 5021 8692 5055
rect 8634 4987 8692 5021
rect 8634 4953 8646 4987
rect 8680 4953 8692 4987
rect 8634 4919 8692 4953
rect 8634 4885 8646 4919
rect 8680 4885 8692 4919
rect 8634 4851 8692 4885
rect 8634 4817 8646 4851
rect 8680 4817 8692 4851
rect 8634 4783 8692 4817
rect 8634 4749 8646 4783
rect 8680 4749 8692 4783
rect 8634 4715 8692 4749
rect 8634 4681 8646 4715
rect 8680 4681 8692 4715
rect 8634 4647 8692 4681
rect 8634 4613 8646 4647
rect 8680 4613 8692 4647
rect 8634 4579 8692 4613
rect 8634 4545 8646 4579
rect 8680 4545 8692 4579
rect 8634 4511 8692 4545
rect 8634 4477 8646 4511
rect 8680 4477 8692 4511
rect 8634 4443 8692 4477
rect 8634 4409 8646 4443
rect 8680 4409 8692 4443
rect 8634 4375 8692 4409
rect 8634 4341 8646 4375
rect 8680 4341 8692 4375
rect 8634 4307 8692 4341
rect 8634 4273 8646 4307
rect 8680 4273 8692 4307
rect 8634 4239 8692 4273
rect 8634 4205 8646 4239
rect 8680 4205 8692 4239
rect 8634 4171 8692 4205
rect 8634 4137 8646 4171
rect 8680 4137 8692 4171
rect 8634 4103 8692 4137
rect 8634 4069 8646 4103
rect 8680 4069 8692 4103
rect 8634 4035 8692 4069
rect 8634 4001 8646 4035
rect 8680 4001 8692 4035
rect 8634 3967 8692 4001
rect 8634 3933 8646 3967
rect 8680 3933 8692 3967
rect 8634 3899 8692 3933
rect 8634 3865 8646 3899
rect 8680 3865 8692 3899
rect 8634 3831 8692 3865
rect 8634 3797 8646 3831
rect 8680 3797 8692 3831
rect 8634 3763 8692 3797
rect 8634 3729 8646 3763
rect 8680 3729 8692 3763
rect 8634 3695 8692 3729
rect 8634 3661 8646 3695
rect 8680 3661 8692 3695
rect 8634 3630 8692 3661
rect 8892 5599 8950 5630
rect 8892 5565 8904 5599
rect 8938 5565 8950 5599
rect 8892 5531 8950 5565
rect 8892 5497 8904 5531
rect 8938 5497 8950 5531
rect 8892 5463 8950 5497
rect 8892 5429 8904 5463
rect 8938 5429 8950 5463
rect 8892 5395 8950 5429
rect 8892 5361 8904 5395
rect 8938 5361 8950 5395
rect 8892 5327 8950 5361
rect 8892 5293 8904 5327
rect 8938 5293 8950 5327
rect 8892 5259 8950 5293
rect 8892 5225 8904 5259
rect 8938 5225 8950 5259
rect 8892 5191 8950 5225
rect 8892 5157 8904 5191
rect 8938 5157 8950 5191
rect 8892 5123 8950 5157
rect 8892 5089 8904 5123
rect 8938 5089 8950 5123
rect 8892 5055 8950 5089
rect 8892 5021 8904 5055
rect 8938 5021 8950 5055
rect 8892 4987 8950 5021
rect 8892 4953 8904 4987
rect 8938 4953 8950 4987
rect 8892 4919 8950 4953
rect 8892 4885 8904 4919
rect 8938 4885 8950 4919
rect 8892 4851 8950 4885
rect 8892 4817 8904 4851
rect 8938 4817 8950 4851
rect 8892 4783 8950 4817
rect 8892 4749 8904 4783
rect 8938 4749 8950 4783
rect 8892 4715 8950 4749
rect 8892 4681 8904 4715
rect 8938 4681 8950 4715
rect 8892 4647 8950 4681
rect 8892 4613 8904 4647
rect 8938 4613 8950 4647
rect 8892 4579 8950 4613
rect 8892 4545 8904 4579
rect 8938 4545 8950 4579
rect 8892 4511 8950 4545
rect 8892 4477 8904 4511
rect 8938 4477 8950 4511
rect 8892 4443 8950 4477
rect 8892 4409 8904 4443
rect 8938 4409 8950 4443
rect 8892 4375 8950 4409
rect 8892 4341 8904 4375
rect 8938 4341 8950 4375
rect 8892 4307 8950 4341
rect 8892 4273 8904 4307
rect 8938 4273 8950 4307
rect 8892 4239 8950 4273
rect 8892 4205 8904 4239
rect 8938 4205 8950 4239
rect 8892 4171 8950 4205
rect 8892 4137 8904 4171
rect 8938 4137 8950 4171
rect 8892 4103 8950 4137
rect 8892 4069 8904 4103
rect 8938 4069 8950 4103
rect 8892 4035 8950 4069
rect 8892 4001 8904 4035
rect 8938 4001 8950 4035
rect 8892 3967 8950 4001
rect 8892 3933 8904 3967
rect 8938 3933 8950 3967
rect 8892 3899 8950 3933
rect 8892 3865 8904 3899
rect 8938 3865 8950 3899
rect 8892 3831 8950 3865
rect 8892 3797 8904 3831
rect 8938 3797 8950 3831
rect 8892 3763 8950 3797
rect 8892 3729 8904 3763
rect 8938 3729 8950 3763
rect 8892 3695 8950 3729
rect 8892 3661 8904 3695
rect 8938 3661 8950 3695
rect 8892 3630 8950 3661
rect 9334 5599 9392 5630
rect 9334 5565 9346 5599
rect 9380 5565 9392 5599
rect 9334 5531 9392 5565
rect 9334 5497 9346 5531
rect 9380 5497 9392 5531
rect 9334 5463 9392 5497
rect 9334 5429 9346 5463
rect 9380 5429 9392 5463
rect 9334 5395 9392 5429
rect 9334 5361 9346 5395
rect 9380 5361 9392 5395
rect 9334 5327 9392 5361
rect 9334 5293 9346 5327
rect 9380 5293 9392 5327
rect 9334 5259 9392 5293
rect 9334 5225 9346 5259
rect 9380 5225 9392 5259
rect 9334 5191 9392 5225
rect 9334 5157 9346 5191
rect 9380 5157 9392 5191
rect 9334 5123 9392 5157
rect 9334 5089 9346 5123
rect 9380 5089 9392 5123
rect 9334 5055 9392 5089
rect 9334 5021 9346 5055
rect 9380 5021 9392 5055
rect 9334 4987 9392 5021
rect 9334 4953 9346 4987
rect 9380 4953 9392 4987
rect 9334 4919 9392 4953
rect 9334 4885 9346 4919
rect 9380 4885 9392 4919
rect 9334 4851 9392 4885
rect 9334 4817 9346 4851
rect 9380 4817 9392 4851
rect 9334 4783 9392 4817
rect 9334 4749 9346 4783
rect 9380 4749 9392 4783
rect 9334 4715 9392 4749
rect 9334 4681 9346 4715
rect 9380 4681 9392 4715
rect 9334 4647 9392 4681
rect 9334 4613 9346 4647
rect 9380 4613 9392 4647
rect 9334 4579 9392 4613
rect 9334 4545 9346 4579
rect 9380 4545 9392 4579
rect 9334 4511 9392 4545
rect 9334 4477 9346 4511
rect 9380 4477 9392 4511
rect 9334 4443 9392 4477
rect 9334 4409 9346 4443
rect 9380 4409 9392 4443
rect 9334 4375 9392 4409
rect 9334 4341 9346 4375
rect 9380 4341 9392 4375
rect 9334 4307 9392 4341
rect 9334 4273 9346 4307
rect 9380 4273 9392 4307
rect 9334 4239 9392 4273
rect 9334 4205 9346 4239
rect 9380 4205 9392 4239
rect 9334 4171 9392 4205
rect 9334 4137 9346 4171
rect 9380 4137 9392 4171
rect 9334 4103 9392 4137
rect 9334 4069 9346 4103
rect 9380 4069 9392 4103
rect 9334 4035 9392 4069
rect 9334 4001 9346 4035
rect 9380 4001 9392 4035
rect 9334 3967 9392 4001
rect 9334 3933 9346 3967
rect 9380 3933 9392 3967
rect 9334 3899 9392 3933
rect 9334 3865 9346 3899
rect 9380 3865 9392 3899
rect 9334 3831 9392 3865
rect 9334 3797 9346 3831
rect 9380 3797 9392 3831
rect 9334 3763 9392 3797
rect 9334 3729 9346 3763
rect 9380 3729 9392 3763
rect 9334 3695 9392 3729
rect 9334 3661 9346 3695
rect 9380 3661 9392 3695
rect 9334 3630 9392 3661
rect 9592 5599 9650 5630
rect 9592 5565 9604 5599
rect 9638 5565 9650 5599
rect 9592 5531 9650 5565
rect 9592 5497 9604 5531
rect 9638 5497 9650 5531
rect 9592 5463 9650 5497
rect 9592 5429 9604 5463
rect 9638 5429 9650 5463
rect 9592 5395 9650 5429
rect 9592 5361 9604 5395
rect 9638 5361 9650 5395
rect 9592 5327 9650 5361
rect 9592 5293 9604 5327
rect 9638 5293 9650 5327
rect 9592 5259 9650 5293
rect 9592 5225 9604 5259
rect 9638 5225 9650 5259
rect 9592 5191 9650 5225
rect 9592 5157 9604 5191
rect 9638 5157 9650 5191
rect 9592 5123 9650 5157
rect 9592 5089 9604 5123
rect 9638 5089 9650 5123
rect 9592 5055 9650 5089
rect 9592 5021 9604 5055
rect 9638 5021 9650 5055
rect 9592 4987 9650 5021
rect 9592 4953 9604 4987
rect 9638 4953 9650 4987
rect 9592 4919 9650 4953
rect 9592 4885 9604 4919
rect 9638 4885 9650 4919
rect 9592 4851 9650 4885
rect 9592 4817 9604 4851
rect 9638 4817 9650 4851
rect 9592 4783 9650 4817
rect 9592 4749 9604 4783
rect 9638 4749 9650 4783
rect 9592 4715 9650 4749
rect 9592 4681 9604 4715
rect 9638 4681 9650 4715
rect 9592 4647 9650 4681
rect 9592 4613 9604 4647
rect 9638 4613 9650 4647
rect 9592 4579 9650 4613
rect 9592 4545 9604 4579
rect 9638 4545 9650 4579
rect 9592 4511 9650 4545
rect 9592 4477 9604 4511
rect 9638 4477 9650 4511
rect 9592 4443 9650 4477
rect 9592 4409 9604 4443
rect 9638 4409 9650 4443
rect 9592 4375 9650 4409
rect 9592 4341 9604 4375
rect 9638 4341 9650 4375
rect 9592 4307 9650 4341
rect 9592 4273 9604 4307
rect 9638 4273 9650 4307
rect 9592 4239 9650 4273
rect 9592 4205 9604 4239
rect 9638 4205 9650 4239
rect 9592 4171 9650 4205
rect 9592 4137 9604 4171
rect 9638 4137 9650 4171
rect 9592 4103 9650 4137
rect 9592 4069 9604 4103
rect 9638 4069 9650 4103
rect 9592 4035 9650 4069
rect 9592 4001 9604 4035
rect 9638 4001 9650 4035
rect 9592 3967 9650 4001
rect 9592 3933 9604 3967
rect 9638 3933 9650 3967
rect 9592 3899 9650 3933
rect 9592 3865 9604 3899
rect 9638 3865 9650 3899
rect 9592 3831 9650 3865
rect 9592 3797 9604 3831
rect 9638 3797 9650 3831
rect 9592 3763 9650 3797
rect 9592 3729 9604 3763
rect 9638 3729 9650 3763
rect 9592 3695 9650 3729
rect 9592 3661 9604 3695
rect 9638 3661 9650 3695
rect 9592 3630 9650 3661
rect 10034 5599 10092 5630
rect 10034 5565 10046 5599
rect 10080 5565 10092 5599
rect 10034 5531 10092 5565
rect 10034 5497 10046 5531
rect 10080 5497 10092 5531
rect 10034 5463 10092 5497
rect 10034 5429 10046 5463
rect 10080 5429 10092 5463
rect 10034 5395 10092 5429
rect 10034 5361 10046 5395
rect 10080 5361 10092 5395
rect 10034 5327 10092 5361
rect 10034 5293 10046 5327
rect 10080 5293 10092 5327
rect 10034 5259 10092 5293
rect 10034 5225 10046 5259
rect 10080 5225 10092 5259
rect 10034 5191 10092 5225
rect 10034 5157 10046 5191
rect 10080 5157 10092 5191
rect 10034 5123 10092 5157
rect 10034 5089 10046 5123
rect 10080 5089 10092 5123
rect 10034 5055 10092 5089
rect 10034 5021 10046 5055
rect 10080 5021 10092 5055
rect 10034 4987 10092 5021
rect 10034 4953 10046 4987
rect 10080 4953 10092 4987
rect 10034 4919 10092 4953
rect 10034 4885 10046 4919
rect 10080 4885 10092 4919
rect 10034 4851 10092 4885
rect 10034 4817 10046 4851
rect 10080 4817 10092 4851
rect 10034 4783 10092 4817
rect 10034 4749 10046 4783
rect 10080 4749 10092 4783
rect 10034 4715 10092 4749
rect 10034 4681 10046 4715
rect 10080 4681 10092 4715
rect 10034 4647 10092 4681
rect 10034 4613 10046 4647
rect 10080 4613 10092 4647
rect 10034 4579 10092 4613
rect 10034 4545 10046 4579
rect 10080 4545 10092 4579
rect 10034 4511 10092 4545
rect 10034 4477 10046 4511
rect 10080 4477 10092 4511
rect 10034 4443 10092 4477
rect 10034 4409 10046 4443
rect 10080 4409 10092 4443
rect 10034 4375 10092 4409
rect 10034 4341 10046 4375
rect 10080 4341 10092 4375
rect 10034 4307 10092 4341
rect 10034 4273 10046 4307
rect 10080 4273 10092 4307
rect 10034 4239 10092 4273
rect 10034 4205 10046 4239
rect 10080 4205 10092 4239
rect 10034 4171 10092 4205
rect 10034 4137 10046 4171
rect 10080 4137 10092 4171
rect 10034 4103 10092 4137
rect 10034 4069 10046 4103
rect 10080 4069 10092 4103
rect 10034 4035 10092 4069
rect 10034 4001 10046 4035
rect 10080 4001 10092 4035
rect 10034 3967 10092 4001
rect 10034 3933 10046 3967
rect 10080 3933 10092 3967
rect 10034 3899 10092 3933
rect 10034 3865 10046 3899
rect 10080 3865 10092 3899
rect 10034 3831 10092 3865
rect 10034 3797 10046 3831
rect 10080 3797 10092 3831
rect 10034 3763 10092 3797
rect 10034 3729 10046 3763
rect 10080 3729 10092 3763
rect 10034 3695 10092 3729
rect 10034 3661 10046 3695
rect 10080 3661 10092 3695
rect 10034 3630 10092 3661
rect 10292 5599 10350 5630
rect 10292 5565 10304 5599
rect 10338 5565 10350 5599
rect 10292 5531 10350 5565
rect 10292 5497 10304 5531
rect 10338 5497 10350 5531
rect 10292 5463 10350 5497
rect 10292 5429 10304 5463
rect 10338 5429 10350 5463
rect 10292 5395 10350 5429
rect 10292 5361 10304 5395
rect 10338 5361 10350 5395
rect 10292 5327 10350 5361
rect 10292 5293 10304 5327
rect 10338 5293 10350 5327
rect 10292 5259 10350 5293
rect 10292 5225 10304 5259
rect 10338 5225 10350 5259
rect 10292 5191 10350 5225
rect 10292 5157 10304 5191
rect 10338 5157 10350 5191
rect 10292 5123 10350 5157
rect 10292 5089 10304 5123
rect 10338 5089 10350 5123
rect 10292 5055 10350 5089
rect 10292 5021 10304 5055
rect 10338 5021 10350 5055
rect 10292 4987 10350 5021
rect 10292 4953 10304 4987
rect 10338 4953 10350 4987
rect 10292 4919 10350 4953
rect 10292 4885 10304 4919
rect 10338 4885 10350 4919
rect 10292 4851 10350 4885
rect 10292 4817 10304 4851
rect 10338 4817 10350 4851
rect 10292 4783 10350 4817
rect 10292 4749 10304 4783
rect 10338 4749 10350 4783
rect 10292 4715 10350 4749
rect 10292 4681 10304 4715
rect 10338 4681 10350 4715
rect 10292 4647 10350 4681
rect 10292 4613 10304 4647
rect 10338 4613 10350 4647
rect 10292 4579 10350 4613
rect 10292 4545 10304 4579
rect 10338 4545 10350 4579
rect 10292 4511 10350 4545
rect 10292 4477 10304 4511
rect 10338 4477 10350 4511
rect 10292 4443 10350 4477
rect 10292 4409 10304 4443
rect 10338 4409 10350 4443
rect 10292 4375 10350 4409
rect 10292 4341 10304 4375
rect 10338 4341 10350 4375
rect 10292 4307 10350 4341
rect 10292 4273 10304 4307
rect 10338 4273 10350 4307
rect 10292 4239 10350 4273
rect 10292 4205 10304 4239
rect 10338 4205 10350 4239
rect 10292 4171 10350 4205
rect 10292 4137 10304 4171
rect 10338 4137 10350 4171
rect 10292 4103 10350 4137
rect 10292 4069 10304 4103
rect 10338 4069 10350 4103
rect 10292 4035 10350 4069
rect 10292 4001 10304 4035
rect 10338 4001 10350 4035
rect 10292 3967 10350 4001
rect 10292 3933 10304 3967
rect 10338 3933 10350 3967
rect 10292 3899 10350 3933
rect 10292 3865 10304 3899
rect 10338 3865 10350 3899
rect 10292 3831 10350 3865
rect 10292 3797 10304 3831
rect 10338 3797 10350 3831
rect 10292 3763 10350 3797
rect 10292 3729 10304 3763
rect 10338 3729 10350 3763
rect 10292 3695 10350 3729
rect 10292 3661 10304 3695
rect 10338 3661 10350 3695
rect 10292 3630 10350 3661
rect 1076 1901 1134 1916
rect 1076 1867 1088 1901
rect 1122 1867 1134 1901
rect 1076 1833 1134 1867
rect 1076 1799 1088 1833
rect 1122 1799 1134 1833
rect 1076 1765 1134 1799
rect 1076 1731 1088 1765
rect 1122 1731 1134 1765
rect 1076 1716 1134 1731
rect 1534 1901 1592 1916
rect 1534 1867 1546 1901
rect 1580 1867 1592 1901
rect 1534 1833 1592 1867
rect 1534 1799 1546 1833
rect 1580 1799 1592 1833
rect 1534 1765 1592 1799
rect 1534 1731 1546 1765
rect 1580 1731 1592 1765
rect 1534 1716 1592 1731
rect 2076 1901 2134 1916
rect 2076 1867 2088 1901
rect 2122 1867 2134 1901
rect 2076 1833 2134 1867
rect 2076 1799 2088 1833
rect 2122 1799 2134 1833
rect 2076 1765 2134 1799
rect 2076 1731 2088 1765
rect 2122 1731 2134 1765
rect 2076 1716 2134 1731
rect 2534 1901 2592 1916
rect 2534 1867 2546 1901
rect 2580 1867 2592 1901
rect 2534 1833 2592 1867
rect 2534 1799 2546 1833
rect 2580 1799 2592 1833
rect 2534 1765 2592 1799
rect 2534 1731 2546 1765
rect 2580 1731 2592 1765
rect 2534 1716 2592 1731
rect 3076 1901 3134 1916
rect 3076 1867 3088 1901
rect 3122 1867 3134 1901
rect 3076 1833 3134 1867
rect 3076 1799 3088 1833
rect 3122 1799 3134 1833
rect 3076 1765 3134 1799
rect 3076 1731 3088 1765
rect 3122 1731 3134 1765
rect 3076 1716 3134 1731
rect 3534 1901 3592 1916
rect 3534 1867 3546 1901
rect 3580 1867 3592 1901
rect 3534 1833 3592 1867
rect 3534 1799 3546 1833
rect 3580 1799 3592 1833
rect 3534 1765 3592 1799
rect 3534 1731 3546 1765
rect 3580 1731 3592 1765
rect 3534 1716 3592 1731
rect 4076 1901 4134 1916
rect 4076 1867 4088 1901
rect 4122 1867 4134 1901
rect 4076 1833 4134 1867
rect 4076 1799 4088 1833
rect 4122 1799 4134 1833
rect 4076 1765 4134 1799
rect 4076 1731 4088 1765
rect 4122 1731 4134 1765
rect 4076 1716 4134 1731
rect 4534 1901 4592 1916
rect 4534 1867 4546 1901
rect 4580 1867 4592 1901
rect 4534 1833 4592 1867
rect 4534 1799 4546 1833
rect 4580 1799 4592 1833
rect 4534 1765 4592 1799
rect 4534 1731 4546 1765
rect 4580 1731 4592 1765
rect 4534 1716 4592 1731
rect 5076 1901 5134 1916
rect 5076 1867 5088 1901
rect 5122 1867 5134 1901
rect 5076 1833 5134 1867
rect 5076 1799 5088 1833
rect 5122 1799 5134 1833
rect 5076 1765 5134 1799
rect 5076 1731 5088 1765
rect 5122 1731 5134 1765
rect 5076 1716 5134 1731
rect 5534 1901 5592 1916
rect 5534 1867 5546 1901
rect 5580 1867 5592 1901
rect 5534 1833 5592 1867
rect 5534 1799 5546 1833
rect 5580 1799 5592 1833
rect 5534 1765 5592 1799
rect 5534 1731 5546 1765
rect 5580 1731 5592 1765
rect 5534 1716 5592 1731
rect 6076 1901 6134 1916
rect 6076 1867 6088 1901
rect 6122 1867 6134 1901
rect 6076 1833 6134 1867
rect 6076 1799 6088 1833
rect 6122 1799 6134 1833
rect 6076 1765 6134 1799
rect 6076 1731 6088 1765
rect 6122 1731 6134 1765
rect 6076 1716 6134 1731
rect 6534 1901 6592 1916
rect 6534 1867 6546 1901
rect 6580 1867 6592 1901
rect 6534 1833 6592 1867
rect 6534 1799 6546 1833
rect 6580 1799 6592 1833
rect 6534 1765 6592 1799
rect 6534 1731 6546 1765
rect 6580 1731 6592 1765
rect 6534 1716 6592 1731
rect 7076 1901 7134 1916
rect 7076 1867 7088 1901
rect 7122 1867 7134 1901
rect 7076 1833 7134 1867
rect 7076 1799 7088 1833
rect 7122 1799 7134 1833
rect 7076 1765 7134 1799
rect 7076 1731 7088 1765
rect 7122 1731 7134 1765
rect 7076 1716 7134 1731
rect 7534 1901 7592 1916
rect 7534 1867 7546 1901
rect 7580 1867 7592 1901
rect 7534 1833 7592 1867
rect 7534 1799 7546 1833
rect 7580 1799 7592 1833
rect 7534 1765 7592 1799
rect 7534 1731 7546 1765
rect 7580 1731 7592 1765
rect 7534 1716 7592 1731
rect 8076 1901 8134 1916
rect 8076 1867 8088 1901
rect 8122 1867 8134 1901
rect 8076 1833 8134 1867
rect 8076 1799 8088 1833
rect 8122 1799 8134 1833
rect 8076 1765 8134 1799
rect 8076 1731 8088 1765
rect 8122 1731 8134 1765
rect 8076 1716 8134 1731
rect 8534 1901 8592 1916
rect 8534 1867 8546 1901
rect 8580 1867 8592 1901
rect 8534 1833 8592 1867
rect 8534 1799 8546 1833
rect 8580 1799 8592 1833
rect 8534 1765 8592 1799
rect 8534 1731 8546 1765
rect 8580 1731 8592 1765
rect 8534 1716 8592 1731
rect 9076 1901 9134 1916
rect 9076 1867 9088 1901
rect 9122 1867 9134 1901
rect 9076 1833 9134 1867
rect 9076 1799 9088 1833
rect 9122 1799 9134 1833
rect 9076 1765 9134 1799
rect 9076 1731 9088 1765
rect 9122 1731 9134 1765
rect 9076 1716 9134 1731
rect 9534 1901 9592 1916
rect 9534 1867 9546 1901
rect 9580 1867 9592 1901
rect 9534 1833 9592 1867
rect 9534 1799 9546 1833
rect 9580 1799 9592 1833
rect 9534 1765 9592 1799
rect 9534 1731 9546 1765
rect 9580 1731 9592 1765
rect 9534 1716 9592 1731
rect 10076 1901 10134 1916
rect 10076 1867 10088 1901
rect 10122 1867 10134 1901
rect 10076 1833 10134 1867
rect 10076 1799 10088 1833
rect 10122 1799 10134 1833
rect 10076 1765 10134 1799
rect 10076 1731 10088 1765
rect 10122 1731 10134 1765
rect 10076 1716 10134 1731
rect 10534 1901 10592 1916
rect 10534 1867 10546 1901
rect 10580 1867 10592 1901
rect 10534 1833 10592 1867
rect 10534 1799 10546 1833
rect 10580 1799 10592 1833
rect 10534 1765 10592 1799
rect 10534 1731 10546 1765
rect 10580 1731 10592 1765
rect 10534 1716 10592 1731
rect 1076 1401 1134 1416
rect 1076 1367 1088 1401
rect 1122 1367 1134 1401
rect 1076 1333 1134 1367
rect 1076 1299 1088 1333
rect 1122 1299 1134 1333
rect 1076 1265 1134 1299
rect 1076 1231 1088 1265
rect 1122 1231 1134 1265
rect 1076 1216 1134 1231
rect 1534 1401 1592 1416
rect 1534 1367 1546 1401
rect 1580 1367 1592 1401
rect 1534 1333 1592 1367
rect 1534 1299 1546 1333
rect 1580 1299 1592 1333
rect 1534 1265 1592 1299
rect 1534 1231 1546 1265
rect 1580 1231 1592 1265
rect 1534 1216 1592 1231
rect 2076 1401 2134 1416
rect 2076 1367 2088 1401
rect 2122 1367 2134 1401
rect 2076 1333 2134 1367
rect 2076 1299 2088 1333
rect 2122 1299 2134 1333
rect 2076 1265 2134 1299
rect 2076 1231 2088 1265
rect 2122 1231 2134 1265
rect 2076 1216 2134 1231
rect 2534 1401 2592 1416
rect 2534 1367 2546 1401
rect 2580 1367 2592 1401
rect 2534 1333 2592 1367
rect 2534 1299 2546 1333
rect 2580 1299 2592 1333
rect 2534 1265 2592 1299
rect 2534 1231 2546 1265
rect 2580 1231 2592 1265
rect 2534 1216 2592 1231
rect 3076 1401 3134 1416
rect 3076 1367 3088 1401
rect 3122 1367 3134 1401
rect 3076 1333 3134 1367
rect 3076 1299 3088 1333
rect 3122 1299 3134 1333
rect 3076 1265 3134 1299
rect 3076 1231 3088 1265
rect 3122 1231 3134 1265
rect 3076 1216 3134 1231
rect 3534 1401 3592 1416
rect 3534 1367 3546 1401
rect 3580 1367 3592 1401
rect 3534 1333 3592 1367
rect 3534 1299 3546 1333
rect 3580 1299 3592 1333
rect 3534 1265 3592 1299
rect 3534 1231 3546 1265
rect 3580 1231 3592 1265
rect 3534 1216 3592 1231
rect 4076 1401 4134 1416
rect 4076 1367 4088 1401
rect 4122 1367 4134 1401
rect 4076 1333 4134 1367
rect 4076 1299 4088 1333
rect 4122 1299 4134 1333
rect 4076 1265 4134 1299
rect 4076 1231 4088 1265
rect 4122 1231 4134 1265
rect 4076 1216 4134 1231
rect 4534 1401 4592 1416
rect 4534 1367 4546 1401
rect 4580 1367 4592 1401
rect 4534 1333 4592 1367
rect 4534 1299 4546 1333
rect 4580 1299 4592 1333
rect 4534 1265 4592 1299
rect 4534 1231 4546 1265
rect 4580 1231 4592 1265
rect 4534 1216 4592 1231
rect 5076 1401 5134 1416
rect 5076 1367 5088 1401
rect 5122 1367 5134 1401
rect 5076 1333 5134 1367
rect 5076 1299 5088 1333
rect 5122 1299 5134 1333
rect 5076 1265 5134 1299
rect 5076 1231 5088 1265
rect 5122 1231 5134 1265
rect 5076 1216 5134 1231
rect 5534 1401 5592 1416
rect 5534 1367 5546 1401
rect 5580 1367 5592 1401
rect 5534 1333 5592 1367
rect 5534 1299 5546 1333
rect 5580 1299 5592 1333
rect 5534 1265 5592 1299
rect 5534 1231 5546 1265
rect 5580 1231 5592 1265
rect 5534 1216 5592 1231
rect 6076 1401 6134 1416
rect 6076 1367 6088 1401
rect 6122 1367 6134 1401
rect 6076 1333 6134 1367
rect 6076 1299 6088 1333
rect 6122 1299 6134 1333
rect 6076 1265 6134 1299
rect 6076 1231 6088 1265
rect 6122 1231 6134 1265
rect 6076 1216 6134 1231
rect 6534 1401 6592 1416
rect 6534 1367 6546 1401
rect 6580 1367 6592 1401
rect 6534 1333 6592 1367
rect 6534 1299 6546 1333
rect 6580 1299 6592 1333
rect 6534 1265 6592 1299
rect 6534 1231 6546 1265
rect 6580 1231 6592 1265
rect 6534 1216 6592 1231
rect 7076 1401 7134 1416
rect 7076 1367 7088 1401
rect 7122 1367 7134 1401
rect 7076 1333 7134 1367
rect 7076 1299 7088 1333
rect 7122 1299 7134 1333
rect 7076 1265 7134 1299
rect 7076 1231 7088 1265
rect 7122 1231 7134 1265
rect 7076 1216 7134 1231
rect 7534 1401 7592 1416
rect 7534 1367 7546 1401
rect 7580 1367 7592 1401
rect 7534 1333 7592 1367
rect 7534 1299 7546 1333
rect 7580 1299 7592 1333
rect 7534 1265 7592 1299
rect 7534 1231 7546 1265
rect 7580 1231 7592 1265
rect 7534 1216 7592 1231
rect 8076 1401 8134 1416
rect 8076 1367 8088 1401
rect 8122 1367 8134 1401
rect 8076 1333 8134 1367
rect 8076 1299 8088 1333
rect 8122 1299 8134 1333
rect 8076 1265 8134 1299
rect 8076 1231 8088 1265
rect 8122 1231 8134 1265
rect 8076 1216 8134 1231
rect 8534 1401 8592 1416
rect 8534 1367 8546 1401
rect 8580 1367 8592 1401
rect 8534 1333 8592 1367
rect 8534 1299 8546 1333
rect 8580 1299 8592 1333
rect 8534 1265 8592 1299
rect 8534 1231 8546 1265
rect 8580 1231 8592 1265
rect 8534 1216 8592 1231
rect 9076 1401 9134 1416
rect 9076 1367 9088 1401
rect 9122 1367 9134 1401
rect 9076 1333 9134 1367
rect 9076 1299 9088 1333
rect 9122 1299 9134 1333
rect 9076 1265 9134 1299
rect 9076 1231 9088 1265
rect 9122 1231 9134 1265
rect 9076 1216 9134 1231
rect 9534 1401 9592 1416
rect 9534 1367 9546 1401
rect 9580 1367 9592 1401
rect 9534 1333 9592 1367
rect 9534 1299 9546 1333
rect 9580 1299 9592 1333
rect 9534 1265 9592 1299
rect 9534 1231 9546 1265
rect 9580 1231 9592 1265
rect 9534 1216 9592 1231
rect 10076 1401 10134 1416
rect 10076 1367 10088 1401
rect 10122 1367 10134 1401
rect 10076 1333 10134 1367
rect 10076 1299 10088 1333
rect 10122 1299 10134 1333
rect 10076 1265 10134 1299
rect 10076 1231 10088 1265
rect 10122 1231 10134 1265
rect 10076 1216 10134 1231
rect 10534 1401 10592 1416
rect 10534 1367 10546 1401
rect 10580 1367 10592 1401
rect 10534 1333 10592 1367
rect 10534 1299 10546 1333
rect 10580 1299 10592 1333
rect 10534 1265 10592 1299
rect 10534 1231 10546 1265
rect 10580 1231 10592 1265
rect 10534 1216 10592 1231
<< mvpdiff >>
rect 1966 8496 2024 8509
rect 1966 8462 1978 8496
rect 2012 8462 2024 8496
rect 1966 8428 2024 8462
rect 1966 8394 1978 8428
rect 2012 8394 2024 8428
rect 1966 8360 2024 8394
rect 1966 8326 1978 8360
rect 2012 8326 2024 8360
rect 1966 8292 2024 8326
rect 1966 8258 1978 8292
rect 2012 8258 2024 8292
rect 1966 8224 2024 8258
rect 1966 8190 1978 8224
rect 2012 8190 2024 8224
rect 1966 8156 2024 8190
rect 1966 8122 1978 8156
rect 2012 8122 2024 8156
rect 1966 8109 2024 8122
rect 2424 8496 2482 8509
rect 2424 8462 2436 8496
rect 2470 8462 2482 8496
rect 2424 8428 2482 8462
rect 2424 8394 2436 8428
rect 2470 8394 2482 8428
rect 2424 8360 2482 8394
rect 2424 8326 2436 8360
rect 2470 8326 2482 8360
rect 2424 8292 2482 8326
rect 2424 8258 2436 8292
rect 2470 8258 2482 8292
rect 2424 8224 2482 8258
rect 2424 8190 2436 8224
rect 2470 8190 2482 8224
rect 2424 8156 2482 8190
rect 2424 8122 2436 8156
rect 2470 8122 2482 8156
rect 2424 8109 2482 8122
rect 2966 8496 3024 8509
rect 2966 8462 2978 8496
rect 3012 8462 3024 8496
rect 2966 8428 3024 8462
rect 2966 8394 2978 8428
rect 3012 8394 3024 8428
rect 2966 8360 3024 8394
rect 2966 8326 2978 8360
rect 3012 8326 3024 8360
rect 2966 8292 3024 8326
rect 2966 8258 2978 8292
rect 3012 8258 3024 8292
rect 2966 8224 3024 8258
rect 2966 8190 2978 8224
rect 3012 8190 3024 8224
rect 2966 8156 3024 8190
rect 2966 8122 2978 8156
rect 3012 8122 3024 8156
rect 2966 8109 3024 8122
rect 3424 8496 3482 8509
rect 3424 8462 3436 8496
rect 3470 8462 3482 8496
rect 3424 8428 3482 8462
rect 3424 8394 3436 8428
rect 3470 8394 3482 8428
rect 3424 8360 3482 8394
rect 3424 8326 3436 8360
rect 3470 8326 3482 8360
rect 3424 8292 3482 8326
rect 3424 8258 3436 8292
rect 3470 8258 3482 8292
rect 3424 8224 3482 8258
rect 3424 8190 3436 8224
rect 3470 8190 3482 8224
rect 3424 8156 3482 8190
rect 3424 8122 3436 8156
rect 3470 8122 3482 8156
rect 3424 8109 3482 8122
rect 1966 7756 2024 7769
rect 1966 7722 1978 7756
rect 2012 7722 2024 7756
rect 1966 7688 2024 7722
rect 1966 7654 1978 7688
rect 2012 7654 2024 7688
rect 1966 7620 2024 7654
rect 1966 7586 1978 7620
rect 2012 7586 2024 7620
rect 1966 7552 2024 7586
rect 1966 7518 1978 7552
rect 2012 7518 2024 7552
rect 1966 7484 2024 7518
rect 1966 7450 1978 7484
rect 2012 7450 2024 7484
rect 1966 7416 2024 7450
rect 1966 7382 1978 7416
rect 2012 7382 2024 7416
rect 1966 7369 2024 7382
rect 2424 7756 2482 7769
rect 2424 7722 2436 7756
rect 2470 7722 2482 7756
rect 2424 7688 2482 7722
rect 2424 7654 2436 7688
rect 2470 7654 2482 7688
rect 2424 7620 2482 7654
rect 2424 7586 2436 7620
rect 2470 7586 2482 7620
rect 2424 7552 2482 7586
rect 2424 7518 2436 7552
rect 2470 7518 2482 7552
rect 2424 7484 2482 7518
rect 2424 7450 2436 7484
rect 2470 7450 2482 7484
rect 2424 7416 2482 7450
rect 2424 7382 2436 7416
rect 2470 7382 2482 7416
rect 2424 7369 2482 7382
rect 2966 7756 3024 7769
rect 2966 7722 2978 7756
rect 3012 7722 3024 7756
rect 2966 7688 3024 7722
rect 2966 7654 2978 7688
rect 3012 7654 3024 7688
rect 2966 7620 3024 7654
rect 2966 7586 2978 7620
rect 3012 7586 3024 7620
rect 2966 7552 3024 7586
rect 2966 7518 2978 7552
rect 3012 7518 3024 7552
rect 2966 7484 3024 7518
rect 2966 7450 2978 7484
rect 3012 7450 3024 7484
rect 2966 7416 3024 7450
rect 2966 7382 2978 7416
rect 3012 7382 3024 7416
rect 2966 7369 3024 7382
rect 3424 7756 3482 7769
rect 3424 7722 3436 7756
rect 3470 7722 3482 7756
rect 3424 7688 3482 7722
rect 3424 7654 3436 7688
rect 3470 7654 3482 7688
rect 3424 7620 3482 7654
rect 3424 7586 3436 7620
rect 3470 7586 3482 7620
rect 3424 7552 3482 7586
rect 3424 7518 3436 7552
rect 3470 7518 3482 7552
rect 3424 7484 3482 7518
rect 3424 7450 3436 7484
rect 3470 7450 3482 7484
rect 3424 7416 3482 7450
rect 3424 7382 3436 7416
rect 3470 7382 3482 7416
rect 3424 7369 3482 7382
rect 11684 6836 11742 6849
rect 11684 6802 11696 6836
rect 11730 6802 11742 6836
rect 11684 6768 11742 6802
rect 11684 6734 11696 6768
rect 11730 6734 11742 6768
rect 11684 6700 11742 6734
rect 11684 6666 11696 6700
rect 11730 6666 11742 6700
rect 11684 6632 11742 6666
rect 11684 6598 11696 6632
rect 11730 6598 11742 6632
rect 11684 6564 11742 6598
rect 11684 6530 11696 6564
rect 11730 6530 11742 6564
rect 11684 6496 11742 6530
rect 11684 6462 11696 6496
rect 11730 6462 11742 6496
rect 11684 6449 11742 6462
rect 12142 6836 12200 6849
rect 12142 6802 12154 6836
rect 12188 6802 12200 6836
rect 12142 6768 12200 6802
rect 12142 6734 12154 6768
rect 12188 6734 12200 6768
rect 12142 6700 12200 6734
rect 12142 6666 12154 6700
rect 12188 6666 12200 6700
rect 12142 6632 12200 6666
rect 12142 6598 12154 6632
rect 12188 6598 12200 6632
rect 12142 6564 12200 6598
rect 12142 6530 12154 6564
rect 12188 6530 12200 6564
rect 12142 6496 12200 6530
rect 12142 6462 12154 6496
rect 12188 6462 12200 6496
rect 12142 6449 12200 6462
rect 12584 6836 12642 6849
rect 12584 6802 12596 6836
rect 12630 6802 12642 6836
rect 12584 6768 12642 6802
rect 12584 6734 12596 6768
rect 12630 6734 12642 6768
rect 12584 6700 12642 6734
rect 12584 6666 12596 6700
rect 12630 6666 12642 6700
rect 12584 6632 12642 6666
rect 12584 6598 12596 6632
rect 12630 6598 12642 6632
rect 12584 6564 12642 6598
rect 12584 6530 12596 6564
rect 12630 6530 12642 6564
rect 12584 6496 12642 6530
rect 12584 6462 12596 6496
rect 12630 6462 12642 6496
rect 12584 6449 12642 6462
rect 13042 6836 13100 6849
rect 13042 6802 13054 6836
rect 13088 6802 13100 6836
rect 13042 6768 13100 6802
rect 13042 6734 13054 6768
rect 13088 6734 13100 6768
rect 13042 6700 13100 6734
rect 13042 6666 13054 6700
rect 13088 6666 13100 6700
rect 13042 6632 13100 6666
rect 13042 6598 13054 6632
rect 13088 6598 13100 6632
rect 13042 6564 13100 6598
rect 13042 6530 13054 6564
rect 13088 6530 13100 6564
rect 13042 6496 13100 6530
rect 13042 6462 13054 6496
rect 13088 6462 13100 6496
rect 13042 6449 13100 6462
rect 13484 6836 13542 6849
rect 13484 6802 13496 6836
rect 13530 6802 13542 6836
rect 13484 6768 13542 6802
rect 13484 6734 13496 6768
rect 13530 6734 13542 6768
rect 13484 6700 13542 6734
rect 13484 6666 13496 6700
rect 13530 6666 13542 6700
rect 13484 6632 13542 6666
rect 13484 6598 13496 6632
rect 13530 6598 13542 6632
rect 13484 6564 13542 6598
rect 13484 6530 13496 6564
rect 13530 6530 13542 6564
rect 13484 6496 13542 6530
rect 13484 6462 13496 6496
rect 13530 6462 13542 6496
rect 13484 6449 13542 6462
rect 13942 6836 14000 6849
rect 13942 6802 13954 6836
rect 13988 6802 14000 6836
rect 13942 6768 14000 6802
rect 13942 6734 13954 6768
rect 13988 6734 14000 6768
rect 13942 6700 14000 6734
rect 13942 6666 13954 6700
rect 13988 6666 14000 6700
rect 13942 6632 14000 6666
rect 13942 6598 13954 6632
rect 13988 6598 14000 6632
rect 13942 6564 14000 6598
rect 13942 6530 13954 6564
rect 13988 6530 14000 6564
rect 13942 6496 14000 6530
rect 13942 6462 13954 6496
rect 13988 6462 14000 6496
rect 13942 6449 14000 6462
rect 14384 6836 14442 6849
rect 14384 6802 14396 6836
rect 14430 6802 14442 6836
rect 14384 6768 14442 6802
rect 14384 6734 14396 6768
rect 14430 6734 14442 6768
rect 14384 6700 14442 6734
rect 14384 6666 14396 6700
rect 14430 6666 14442 6700
rect 14384 6632 14442 6666
rect 14384 6598 14396 6632
rect 14430 6598 14442 6632
rect 14384 6564 14442 6598
rect 14384 6530 14396 6564
rect 14430 6530 14442 6564
rect 14384 6496 14442 6530
rect 14384 6462 14396 6496
rect 14430 6462 14442 6496
rect 14384 6449 14442 6462
rect 14842 6836 14900 6849
rect 14842 6802 14854 6836
rect 14888 6802 14900 6836
rect 14842 6768 14900 6802
rect 14842 6734 14854 6768
rect 14888 6734 14900 6768
rect 14842 6700 14900 6734
rect 14842 6666 14854 6700
rect 14888 6666 14900 6700
rect 14842 6632 14900 6666
rect 14842 6598 14854 6632
rect 14888 6598 14900 6632
rect 14842 6564 14900 6598
rect 14842 6530 14854 6564
rect 14888 6530 14900 6564
rect 14842 6496 14900 6530
rect 14842 6462 14854 6496
rect 14888 6462 14900 6496
rect 14842 6449 14900 6462
rect 15284 6836 15342 6849
rect 15284 6802 15296 6836
rect 15330 6802 15342 6836
rect 15284 6768 15342 6802
rect 15284 6734 15296 6768
rect 15330 6734 15342 6768
rect 15284 6700 15342 6734
rect 15284 6666 15296 6700
rect 15330 6666 15342 6700
rect 15284 6632 15342 6666
rect 15284 6598 15296 6632
rect 15330 6598 15342 6632
rect 15284 6564 15342 6598
rect 15284 6530 15296 6564
rect 15330 6530 15342 6564
rect 15284 6496 15342 6530
rect 15284 6462 15296 6496
rect 15330 6462 15342 6496
rect 15284 6449 15342 6462
rect 15742 6836 15800 6849
rect 15742 6802 15754 6836
rect 15788 6802 15800 6836
rect 15742 6768 15800 6802
rect 15742 6734 15754 6768
rect 15788 6734 15800 6768
rect 15742 6700 15800 6734
rect 15742 6666 15754 6700
rect 15788 6666 15800 6700
rect 15742 6632 15800 6666
rect 15742 6598 15754 6632
rect 15788 6598 15800 6632
rect 15742 6564 15800 6598
rect 15742 6530 15754 6564
rect 15788 6530 15800 6564
rect 15742 6496 15800 6530
rect 15742 6462 15754 6496
rect 15788 6462 15800 6496
rect 15742 6449 15800 6462
rect 16184 6836 16242 6849
rect 16184 6802 16196 6836
rect 16230 6802 16242 6836
rect 16184 6768 16242 6802
rect 16184 6734 16196 6768
rect 16230 6734 16242 6768
rect 16184 6700 16242 6734
rect 16184 6666 16196 6700
rect 16230 6666 16242 6700
rect 16184 6632 16242 6666
rect 16184 6598 16196 6632
rect 16230 6598 16242 6632
rect 16184 6564 16242 6598
rect 16184 6530 16196 6564
rect 16230 6530 16242 6564
rect 16184 6496 16242 6530
rect 16184 6462 16196 6496
rect 16230 6462 16242 6496
rect 16184 6449 16242 6462
rect 16642 6836 16700 6849
rect 16642 6802 16654 6836
rect 16688 6802 16700 6836
rect 16642 6768 16700 6802
rect 16642 6734 16654 6768
rect 16688 6734 16700 6768
rect 16642 6700 16700 6734
rect 16642 6666 16654 6700
rect 16688 6666 16700 6700
rect 16642 6632 16700 6666
rect 16642 6598 16654 6632
rect 16688 6598 16700 6632
rect 16642 6564 16700 6598
rect 16642 6530 16654 6564
rect 16688 6530 16700 6564
rect 16642 6496 16700 6530
rect 16642 6462 16654 6496
rect 16688 6462 16700 6496
rect 16642 6449 16700 6462
rect 17084 6836 17142 6849
rect 17084 6802 17096 6836
rect 17130 6802 17142 6836
rect 17084 6768 17142 6802
rect 17084 6734 17096 6768
rect 17130 6734 17142 6768
rect 17084 6700 17142 6734
rect 17084 6666 17096 6700
rect 17130 6666 17142 6700
rect 17084 6632 17142 6666
rect 17084 6598 17096 6632
rect 17130 6598 17142 6632
rect 17084 6564 17142 6598
rect 17084 6530 17096 6564
rect 17130 6530 17142 6564
rect 17084 6496 17142 6530
rect 17084 6462 17096 6496
rect 17130 6462 17142 6496
rect 17084 6449 17142 6462
rect 17542 6836 17600 6849
rect 17542 6802 17554 6836
rect 17588 6802 17600 6836
rect 17542 6768 17600 6802
rect 17542 6734 17554 6768
rect 17588 6734 17600 6768
rect 17542 6700 17600 6734
rect 17542 6666 17554 6700
rect 17588 6666 17600 6700
rect 17542 6632 17600 6666
rect 17542 6598 17554 6632
rect 17588 6598 17600 6632
rect 17542 6564 17600 6598
rect 17542 6530 17554 6564
rect 17588 6530 17600 6564
rect 17542 6496 17600 6530
rect 17542 6462 17554 6496
rect 17588 6462 17600 6496
rect 17542 6449 17600 6462
rect 17984 6836 18042 6849
rect 17984 6802 17996 6836
rect 18030 6802 18042 6836
rect 17984 6768 18042 6802
rect 17984 6734 17996 6768
rect 18030 6734 18042 6768
rect 17984 6700 18042 6734
rect 17984 6666 17996 6700
rect 18030 6666 18042 6700
rect 17984 6632 18042 6666
rect 17984 6598 17996 6632
rect 18030 6598 18042 6632
rect 17984 6564 18042 6598
rect 17984 6530 17996 6564
rect 18030 6530 18042 6564
rect 17984 6496 18042 6530
rect 17984 6462 17996 6496
rect 18030 6462 18042 6496
rect 17984 6449 18042 6462
rect 18442 6836 18500 6849
rect 18442 6802 18454 6836
rect 18488 6802 18500 6836
rect 18442 6768 18500 6802
rect 18442 6734 18454 6768
rect 18488 6734 18500 6768
rect 18442 6700 18500 6734
rect 18442 6666 18454 6700
rect 18488 6666 18500 6700
rect 18442 6632 18500 6666
rect 18442 6598 18454 6632
rect 18488 6598 18500 6632
rect 18442 6564 18500 6598
rect 18442 6530 18454 6564
rect 18488 6530 18500 6564
rect 18442 6496 18500 6530
rect 18442 6462 18454 6496
rect 18488 6462 18500 6496
rect 18442 6449 18500 6462
rect 11684 6096 11742 6109
rect 11684 6062 11696 6096
rect 11730 6062 11742 6096
rect 11684 6028 11742 6062
rect 11684 5994 11696 6028
rect 11730 5994 11742 6028
rect 11684 5960 11742 5994
rect 11684 5926 11696 5960
rect 11730 5926 11742 5960
rect 11684 5892 11742 5926
rect 11684 5858 11696 5892
rect 11730 5858 11742 5892
rect 11684 5824 11742 5858
rect 11684 5790 11696 5824
rect 11730 5790 11742 5824
rect 11684 5756 11742 5790
rect 11684 5722 11696 5756
rect 11730 5722 11742 5756
rect 11684 5709 11742 5722
rect 12142 6096 12200 6109
rect 12142 6062 12154 6096
rect 12188 6062 12200 6096
rect 12142 6028 12200 6062
rect 12142 5994 12154 6028
rect 12188 5994 12200 6028
rect 12142 5960 12200 5994
rect 12142 5926 12154 5960
rect 12188 5926 12200 5960
rect 12142 5892 12200 5926
rect 12142 5858 12154 5892
rect 12188 5858 12200 5892
rect 12142 5824 12200 5858
rect 12142 5790 12154 5824
rect 12188 5790 12200 5824
rect 12142 5756 12200 5790
rect 12142 5722 12154 5756
rect 12188 5722 12200 5756
rect 12142 5709 12200 5722
rect 12584 6096 12642 6109
rect 12584 6062 12596 6096
rect 12630 6062 12642 6096
rect 12584 6028 12642 6062
rect 12584 5994 12596 6028
rect 12630 5994 12642 6028
rect 12584 5960 12642 5994
rect 12584 5926 12596 5960
rect 12630 5926 12642 5960
rect 12584 5892 12642 5926
rect 12584 5858 12596 5892
rect 12630 5858 12642 5892
rect 12584 5824 12642 5858
rect 12584 5790 12596 5824
rect 12630 5790 12642 5824
rect 12584 5756 12642 5790
rect 12584 5722 12596 5756
rect 12630 5722 12642 5756
rect 12584 5709 12642 5722
rect 13042 6096 13100 6109
rect 13042 6062 13054 6096
rect 13088 6062 13100 6096
rect 13042 6028 13100 6062
rect 13042 5994 13054 6028
rect 13088 5994 13100 6028
rect 13042 5960 13100 5994
rect 13042 5926 13054 5960
rect 13088 5926 13100 5960
rect 13042 5892 13100 5926
rect 13042 5858 13054 5892
rect 13088 5858 13100 5892
rect 13042 5824 13100 5858
rect 13042 5790 13054 5824
rect 13088 5790 13100 5824
rect 13042 5756 13100 5790
rect 13042 5722 13054 5756
rect 13088 5722 13100 5756
rect 13042 5709 13100 5722
rect 13484 6096 13542 6109
rect 13484 6062 13496 6096
rect 13530 6062 13542 6096
rect 13484 6028 13542 6062
rect 13484 5994 13496 6028
rect 13530 5994 13542 6028
rect 13484 5960 13542 5994
rect 13484 5926 13496 5960
rect 13530 5926 13542 5960
rect 13484 5892 13542 5926
rect 13484 5858 13496 5892
rect 13530 5858 13542 5892
rect 13484 5824 13542 5858
rect 13484 5790 13496 5824
rect 13530 5790 13542 5824
rect 13484 5756 13542 5790
rect 13484 5722 13496 5756
rect 13530 5722 13542 5756
rect 13484 5709 13542 5722
rect 13942 6096 14000 6109
rect 13942 6062 13954 6096
rect 13988 6062 14000 6096
rect 13942 6028 14000 6062
rect 13942 5994 13954 6028
rect 13988 5994 14000 6028
rect 13942 5960 14000 5994
rect 13942 5926 13954 5960
rect 13988 5926 14000 5960
rect 13942 5892 14000 5926
rect 13942 5858 13954 5892
rect 13988 5858 14000 5892
rect 13942 5824 14000 5858
rect 13942 5790 13954 5824
rect 13988 5790 14000 5824
rect 13942 5756 14000 5790
rect 13942 5722 13954 5756
rect 13988 5722 14000 5756
rect 13942 5709 14000 5722
rect 14384 6096 14442 6109
rect 14384 6062 14396 6096
rect 14430 6062 14442 6096
rect 14384 6028 14442 6062
rect 14384 5994 14396 6028
rect 14430 5994 14442 6028
rect 14384 5960 14442 5994
rect 14384 5926 14396 5960
rect 14430 5926 14442 5960
rect 14384 5892 14442 5926
rect 14384 5858 14396 5892
rect 14430 5858 14442 5892
rect 14384 5824 14442 5858
rect 14384 5790 14396 5824
rect 14430 5790 14442 5824
rect 14384 5756 14442 5790
rect 14384 5722 14396 5756
rect 14430 5722 14442 5756
rect 14384 5709 14442 5722
rect 14842 6096 14900 6109
rect 14842 6062 14854 6096
rect 14888 6062 14900 6096
rect 14842 6028 14900 6062
rect 14842 5994 14854 6028
rect 14888 5994 14900 6028
rect 14842 5960 14900 5994
rect 14842 5926 14854 5960
rect 14888 5926 14900 5960
rect 14842 5892 14900 5926
rect 14842 5858 14854 5892
rect 14888 5858 14900 5892
rect 14842 5824 14900 5858
rect 14842 5790 14854 5824
rect 14888 5790 14900 5824
rect 14842 5756 14900 5790
rect 14842 5722 14854 5756
rect 14888 5722 14900 5756
rect 14842 5709 14900 5722
rect 15284 6096 15342 6109
rect 15284 6062 15296 6096
rect 15330 6062 15342 6096
rect 15284 6028 15342 6062
rect 15284 5994 15296 6028
rect 15330 5994 15342 6028
rect 15284 5960 15342 5994
rect 15284 5926 15296 5960
rect 15330 5926 15342 5960
rect 15284 5892 15342 5926
rect 15284 5858 15296 5892
rect 15330 5858 15342 5892
rect 15284 5824 15342 5858
rect 15284 5790 15296 5824
rect 15330 5790 15342 5824
rect 15284 5756 15342 5790
rect 15284 5722 15296 5756
rect 15330 5722 15342 5756
rect 15284 5709 15342 5722
rect 15742 6096 15800 6109
rect 15742 6062 15754 6096
rect 15788 6062 15800 6096
rect 15742 6028 15800 6062
rect 15742 5994 15754 6028
rect 15788 5994 15800 6028
rect 15742 5960 15800 5994
rect 15742 5926 15754 5960
rect 15788 5926 15800 5960
rect 15742 5892 15800 5926
rect 15742 5858 15754 5892
rect 15788 5858 15800 5892
rect 15742 5824 15800 5858
rect 15742 5790 15754 5824
rect 15788 5790 15800 5824
rect 15742 5756 15800 5790
rect 15742 5722 15754 5756
rect 15788 5722 15800 5756
rect 15742 5709 15800 5722
rect 16184 6096 16242 6109
rect 16184 6062 16196 6096
rect 16230 6062 16242 6096
rect 16184 6028 16242 6062
rect 16184 5994 16196 6028
rect 16230 5994 16242 6028
rect 16184 5960 16242 5994
rect 16184 5926 16196 5960
rect 16230 5926 16242 5960
rect 16184 5892 16242 5926
rect 16184 5858 16196 5892
rect 16230 5858 16242 5892
rect 16184 5824 16242 5858
rect 16184 5790 16196 5824
rect 16230 5790 16242 5824
rect 16184 5756 16242 5790
rect 16184 5722 16196 5756
rect 16230 5722 16242 5756
rect 16184 5709 16242 5722
rect 16642 6096 16700 6109
rect 16642 6062 16654 6096
rect 16688 6062 16700 6096
rect 16642 6028 16700 6062
rect 16642 5994 16654 6028
rect 16688 5994 16700 6028
rect 16642 5960 16700 5994
rect 16642 5926 16654 5960
rect 16688 5926 16700 5960
rect 16642 5892 16700 5926
rect 16642 5858 16654 5892
rect 16688 5858 16700 5892
rect 16642 5824 16700 5858
rect 16642 5790 16654 5824
rect 16688 5790 16700 5824
rect 16642 5756 16700 5790
rect 16642 5722 16654 5756
rect 16688 5722 16700 5756
rect 16642 5709 16700 5722
rect 17084 6096 17142 6109
rect 17084 6062 17096 6096
rect 17130 6062 17142 6096
rect 17084 6028 17142 6062
rect 17084 5994 17096 6028
rect 17130 5994 17142 6028
rect 17084 5960 17142 5994
rect 17084 5926 17096 5960
rect 17130 5926 17142 5960
rect 17084 5892 17142 5926
rect 17084 5858 17096 5892
rect 17130 5858 17142 5892
rect 17084 5824 17142 5858
rect 17084 5790 17096 5824
rect 17130 5790 17142 5824
rect 17084 5756 17142 5790
rect 17084 5722 17096 5756
rect 17130 5722 17142 5756
rect 17084 5709 17142 5722
rect 17542 6096 17600 6109
rect 17542 6062 17554 6096
rect 17588 6062 17600 6096
rect 17542 6028 17600 6062
rect 17542 5994 17554 6028
rect 17588 5994 17600 6028
rect 17542 5960 17600 5994
rect 17542 5926 17554 5960
rect 17588 5926 17600 5960
rect 17542 5892 17600 5926
rect 17542 5858 17554 5892
rect 17588 5858 17600 5892
rect 17542 5824 17600 5858
rect 17542 5790 17554 5824
rect 17588 5790 17600 5824
rect 17542 5756 17600 5790
rect 17542 5722 17554 5756
rect 17588 5722 17600 5756
rect 17542 5709 17600 5722
rect 17984 6096 18042 6109
rect 17984 6062 17996 6096
rect 18030 6062 18042 6096
rect 17984 6028 18042 6062
rect 17984 5994 17996 6028
rect 18030 5994 18042 6028
rect 17984 5960 18042 5994
rect 17984 5926 17996 5960
rect 18030 5926 18042 5960
rect 17984 5892 18042 5926
rect 17984 5858 17996 5892
rect 18030 5858 18042 5892
rect 17984 5824 18042 5858
rect 17984 5790 17996 5824
rect 18030 5790 18042 5824
rect 17984 5756 18042 5790
rect 17984 5722 17996 5756
rect 18030 5722 18042 5756
rect 17984 5709 18042 5722
rect 18442 6096 18500 6109
rect 18442 6062 18454 6096
rect 18488 6062 18500 6096
rect 18442 6028 18500 6062
rect 18442 5994 18454 6028
rect 18488 5994 18500 6028
rect 18442 5960 18500 5994
rect 18442 5926 18454 5960
rect 18488 5926 18500 5960
rect 18442 5892 18500 5926
rect 18442 5858 18454 5892
rect 18488 5858 18500 5892
rect 18442 5824 18500 5858
rect 18442 5790 18454 5824
rect 18488 5790 18500 5824
rect 18442 5756 18500 5790
rect 18442 5722 18454 5756
rect 18488 5722 18500 5756
rect 18442 5709 18500 5722
<< mvndiffc >>
rect -4254 5565 -4220 5599
rect -4254 5497 -4220 5531
rect -4254 5429 -4220 5463
rect -4254 5361 -4220 5395
rect -4254 5293 -4220 5327
rect -4254 5225 -4220 5259
rect -4254 5157 -4220 5191
rect -4254 5089 -4220 5123
rect -4254 5021 -4220 5055
rect -4254 4953 -4220 4987
rect -4254 4885 -4220 4919
rect -4254 4817 -4220 4851
rect -4254 4749 -4220 4783
rect -4254 4681 -4220 4715
rect -4254 4613 -4220 4647
rect -4254 4545 -4220 4579
rect -4254 4477 -4220 4511
rect -4254 4409 -4220 4443
rect -4254 4341 -4220 4375
rect -4254 4273 -4220 4307
rect -4254 4205 -4220 4239
rect -4254 4137 -4220 4171
rect -4254 4069 -4220 4103
rect -4254 4001 -4220 4035
rect -4254 3933 -4220 3967
rect -4254 3865 -4220 3899
rect -4254 3797 -4220 3831
rect -4254 3729 -4220 3763
rect -4254 3661 -4220 3695
rect -3996 5565 -3962 5599
rect -3996 5497 -3962 5531
rect -3996 5429 -3962 5463
rect -3996 5361 -3962 5395
rect -3996 5293 -3962 5327
rect -3996 5225 -3962 5259
rect -3996 5157 -3962 5191
rect -3996 5089 -3962 5123
rect -3996 5021 -3962 5055
rect -3996 4953 -3962 4987
rect -3996 4885 -3962 4919
rect -3996 4817 -3962 4851
rect -3996 4749 -3962 4783
rect -3996 4681 -3962 4715
rect -3996 4613 -3962 4647
rect -3996 4545 -3962 4579
rect -3996 4477 -3962 4511
rect -3996 4409 -3962 4443
rect -3996 4341 -3962 4375
rect -3996 4273 -3962 4307
rect -3996 4205 -3962 4239
rect -3996 4137 -3962 4171
rect -3996 4069 -3962 4103
rect -3996 4001 -3962 4035
rect -3996 3933 -3962 3967
rect -3996 3865 -3962 3899
rect -3996 3797 -3962 3831
rect -3996 3729 -3962 3763
rect -3996 3661 -3962 3695
rect -3554 5565 -3520 5599
rect -3554 5497 -3520 5531
rect -3554 5429 -3520 5463
rect -3554 5361 -3520 5395
rect -3554 5293 -3520 5327
rect -3554 5225 -3520 5259
rect -3554 5157 -3520 5191
rect -3554 5089 -3520 5123
rect -3554 5021 -3520 5055
rect -3554 4953 -3520 4987
rect -3554 4885 -3520 4919
rect -3554 4817 -3520 4851
rect -3554 4749 -3520 4783
rect -3554 4681 -3520 4715
rect -3554 4613 -3520 4647
rect -3554 4545 -3520 4579
rect -3554 4477 -3520 4511
rect -3554 4409 -3520 4443
rect -3554 4341 -3520 4375
rect -3554 4273 -3520 4307
rect -3554 4205 -3520 4239
rect -3554 4137 -3520 4171
rect -3554 4069 -3520 4103
rect -3554 4001 -3520 4035
rect -3554 3933 -3520 3967
rect -3554 3865 -3520 3899
rect -3554 3797 -3520 3831
rect -3554 3729 -3520 3763
rect -3554 3661 -3520 3695
rect -3296 5565 -3262 5599
rect -3296 5497 -3262 5531
rect -3296 5429 -3262 5463
rect -3296 5361 -3262 5395
rect -3296 5293 -3262 5327
rect -3296 5225 -3262 5259
rect -3296 5157 -3262 5191
rect -3296 5089 -3262 5123
rect -3296 5021 -3262 5055
rect -3296 4953 -3262 4987
rect -3296 4885 -3262 4919
rect -3296 4817 -3262 4851
rect -3296 4749 -3262 4783
rect -3296 4681 -3262 4715
rect -3296 4613 -3262 4647
rect -3296 4545 -3262 4579
rect -3296 4477 -3262 4511
rect -3296 4409 -3262 4443
rect -3296 4341 -3262 4375
rect -3296 4273 -3262 4307
rect -3296 4205 -3262 4239
rect -3296 4137 -3262 4171
rect -3296 4069 -3262 4103
rect -3296 4001 -3262 4035
rect -3296 3933 -3262 3967
rect -3296 3865 -3262 3899
rect -3296 3797 -3262 3831
rect -3296 3729 -3262 3763
rect -3296 3661 -3262 3695
rect -2854 5565 -2820 5599
rect -2854 5497 -2820 5531
rect -2854 5429 -2820 5463
rect -2854 5361 -2820 5395
rect -2854 5293 -2820 5327
rect -2854 5225 -2820 5259
rect -2854 5157 -2820 5191
rect -2854 5089 -2820 5123
rect -2854 5021 -2820 5055
rect -2854 4953 -2820 4987
rect -2854 4885 -2820 4919
rect -2854 4817 -2820 4851
rect -2854 4749 -2820 4783
rect -2854 4681 -2820 4715
rect -2854 4613 -2820 4647
rect -2854 4545 -2820 4579
rect -2854 4477 -2820 4511
rect -2854 4409 -2820 4443
rect -2854 4341 -2820 4375
rect -2854 4273 -2820 4307
rect -2854 4205 -2820 4239
rect -2854 4137 -2820 4171
rect -2854 4069 -2820 4103
rect -2854 4001 -2820 4035
rect -2854 3933 -2820 3967
rect -2854 3865 -2820 3899
rect -2854 3797 -2820 3831
rect -2854 3729 -2820 3763
rect -2854 3661 -2820 3695
rect -2596 5565 -2562 5599
rect -2596 5497 -2562 5531
rect -2596 5429 -2562 5463
rect -2596 5361 -2562 5395
rect -2596 5293 -2562 5327
rect -2596 5225 -2562 5259
rect -2596 5157 -2562 5191
rect -2596 5089 -2562 5123
rect -2596 5021 -2562 5055
rect -2596 4953 -2562 4987
rect -2596 4885 -2562 4919
rect -2596 4817 -2562 4851
rect -2596 4749 -2562 4783
rect -2596 4681 -2562 4715
rect -2596 4613 -2562 4647
rect -2596 4545 -2562 4579
rect -2596 4477 -2562 4511
rect -2596 4409 -2562 4443
rect -2596 4341 -2562 4375
rect -2596 4273 -2562 4307
rect -2596 4205 -2562 4239
rect -2596 4137 -2562 4171
rect -2596 4069 -2562 4103
rect -2596 4001 -2562 4035
rect -2596 3933 -2562 3967
rect -2596 3865 -2562 3899
rect -2596 3797 -2562 3831
rect -2596 3729 -2562 3763
rect -2596 3661 -2562 3695
rect -2154 5565 -2120 5599
rect -2154 5497 -2120 5531
rect -2154 5429 -2120 5463
rect -2154 5361 -2120 5395
rect -2154 5293 -2120 5327
rect -2154 5225 -2120 5259
rect -2154 5157 -2120 5191
rect -2154 5089 -2120 5123
rect -2154 5021 -2120 5055
rect -2154 4953 -2120 4987
rect -2154 4885 -2120 4919
rect -2154 4817 -2120 4851
rect -2154 4749 -2120 4783
rect -2154 4681 -2120 4715
rect -2154 4613 -2120 4647
rect -2154 4545 -2120 4579
rect -2154 4477 -2120 4511
rect -2154 4409 -2120 4443
rect -2154 4341 -2120 4375
rect -2154 4273 -2120 4307
rect -2154 4205 -2120 4239
rect -2154 4137 -2120 4171
rect -2154 4069 -2120 4103
rect -2154 4001 -2120 4035
rect -2154 3933 -2120 3967
rect -2154 3865 -2120 3899
rect -2154 3797 -2120 3831
rect -2154 3729 -2120 3763
rect -2154 3661 -2120 3695
rect -1896 5565 -1862 5599
rect -1896 5497 -1862 5531
rect -1896 5429 -1862 5463
rect -1896 5361 -1862 5395
rect -1896 5293 -1862 5327
rect -1896 5225 -1862 5259
rect -1896 5157 -1862 5191
rect -1896 5089 -1862 5123
rect -1896 5021 -1862 5055
rect -1896 4953 -1862 4987
rect -1896 4885 -1862 4919
rect -1896 4817 -1862 4851
rect -1896 4749 -1862 4783
rect -1896 4681 -1862 4715
rect -1896 4613 -1862 4647
rect -1896 4545 -1862 4579
rect -1896 4477 -1862 4511
rect -1896 4409 -1862 4443
rect -1896 4341 -1862 4375
rect -1896 4273 -1862 4307
rect -1896 4205 -1862 4239
rect -1896 4137 -1862 4171
rect -1896 4069 -1862 4103
rect -1896 4001 -1862 4035
rect -1896 3933 -1862 3967
rect -1896 3865 -1862 3899
rect -1896 3797 -1862 3831
rect -1896 3729 -1862 3763
rect -1896 3661 -1862 3695
rect -1454 5565 -1420 5599
rect -1454 5497 -1420 5531
rect -1454 5429 -1420 5463
rect -1454 5361 -1420 5395
rect -1454 5293 -1420 5327
rect -1454 5225 -1420 5259
rect -1454 5157 -1420 5191
rect -1454 5089 -1420 5123
rect -1454 5021 -1420 5055
rect -1454 4953 -1420 4987
rect -1454 4885 -1420 4919
rect -1454 4817 -1420 4851
rect -1454 4749 -1420 4783
rect -1454 4681 -1420 4715
rect -1454 4613 -1420 4647
rect -1454 4545 -1420 4579
rect -1454 4477 -1420 4511
rect -1454 4409 -1420 4443
rect -1454 4341 -1420 4375
rect -1454 4273 -1420 4307
rect -1454 4205 -1420 4239
rect -1454 4137 -1420 4171
rect -1454 4069 -1420 4103
rect -1454 4001 -1420 4035
rect -1454 3933 -1420 3967
rect -1454 3865 -1420 3899
rect -1454 3797 -1420 3831
rect -1454 3729 -1420 3763
rect -1454 3661 -1420 3695
rect -1196 5565 -1162 5599
rect -1196 5497 -1162 5531
rect -1196 5429 -1162 5463
rect -1196 5361 -1162 5395
rect -1196 5293 -1162 5327
rect -1196 5225 -1162 5259
rect -1196 5157 -1162 5191
rect -1196 5089 -1162 5123
rect -1196 5021 -1162 5055
rect -1196 4953 -1162 4987
rect -1196 4885 -1162 4919
rect -1196 4817 -1162 4851
rect -1196 4749 -1162 4783
rect -1196 4681 -1162 4715
rect -1196 4613 -1162 4647
rect -1196 4545 -1162 4579
rect -1196 4477 -1162 4511
rect -1196 4409 -1162 4443
rect -1196 4341 -1162 4375
rect -1196 4273 -1162 4307
rect -1196 4205 -1162 4239
rect -1196 4137 -1162 4171
rect -1196 4069 -1162 4103
rect -1196 4001 -1162 4035
rect -1196 3933 -1162 3967
rect -1196 3865 -1162 3899
rect -1196 3797 -1162 3831
rect -1196 3729 -1162 3763
rect -1196 3661 -1162 3695
rect -754 5565 -720 5599
rect -754 5497 -720 5531
rect -754 5429 -720 5463
rect -754 5361 -720 5395
rect -754 5293 -720 5327
rect -754 5225 -720 5259
rect -754 5157 -720 5191
rect -754 5089 -720 5123
rect -754 5021 -720 5055
rect -754 4953 -720 4987
rect -754 4885 -720 4919
rect -754 4817 -720 4851
rect -754 4749 -720 4783
rect -754 4681 -720 4715
rect -754 4613 -720 4647
rect -754 4545 -720 4579
rect -754 4477 -720 4511
rect -754 4409 -720 4443
rect -754 4341 -720 4375
rect -754 4273 -720 4307
rect -754 4205 -720 4239
rect -754 4137 -720 4171
rect -754 4069 -720 4103
rect -754 4001 -720 4035
rect -754 3933 -720 3967
rect -754 3865 -720 3899
rect -754 3797 -720 3831
rect -754 3729 -720 3763
rect -754 3661 -720 3695
rect -496 5565 -462 5599
rect -496 5497 -462 5531
rect -496 5429 -462 5463
rect -496 5361 -462 5395
rect -496 5293 -462 5327
rect -496 5225 -462 5259
rect -496 5157 -462 5191
rect -496 5089 -462 5123
rect -496 5021 -462 5055
rect -496 4953 -462 4987
rect -496 4885 -462 4919
rect -496 4817 -462 4851
rect -496 4749 -462 4783
rect -496 4681 -462 4715
rect -496 4613 -462 4647
rect -496 4545 -462 4579
rect -496 4477 -462 4511
rect -496 4409 -462 4443
rect -496 4341 -462 4375
rect -496 4273 -462 4307
rect -496 4205 -462 4239
rect -496 4137 -462 4171
rect -496 4069 -462 4103
rect -496 4001 -462 4035
rect -496 3933 -462 3967
rect -496 3865 -462 3899
rect -496 3797 -462 3831
rect -496 3729 -462 3763
rect -496 3661 -462 3695
rect -54 5565 -20 5599
rect -54 5497 -20 5531
rect -54 5429 -20 5463
rect -54 5361 -20 5395
rect -54 5293 -20 5327
rect -54 5225 -20 5259
rect -54 5157 -20 5191
rect -54 5089 -20 5123
rect -54 5021 -20 5055
rect -54 4953 -20 4987
rect -54 4885 -20 4919
rect -54 4817 -20 4851
rect -54 4749 -20 4783
rect -54 4681 -20 4715
rect -54 4613 -20 4647
rect -54 4545 -20 4579
rect -54 4477 -20 4511
rect -54 4409 -20 4443
rect -54 4341 -20 4375
rect -54 4273 -20 4307
rect -54 4205 -20 4239
rect -54 4137 -20 4171
rect -54 4069 -20 4103
rect -54 4001 -20 4035
rect -54 3933 -20 3967
rect -54 3865 -20 3899
rect -54 3797 -20 3831
rect -54 3729 -20 3763
rect -54 3661 -20 3695
rect 204 5565 238 5599
rect 204 5497 238 5531
rect 204 5429 238 5463
rect 204 5361 238 5395
rect 204 5293 238 5327
rect 204 5225 238 5259
rect 204 5157 238 5191
rect 204 5089 238 5123
rect 204 5021 238 5055
rect 204 4953 238 4987
rect 204 4885 238 4919
rect 204 4817 238 4851
rect 204 4749 238 4783
rect 204 4681 238 4715
rect 204 4613 238 4647
rect 204 4545 238 4579
rect 204 4477 238 4511
rect 204 4409 238 4443
rect 204 4341 238 4375
rect 204 4273 238 4307
rect 204 4205 238 4239
rect 204 4137 238 4171
rect 204 4069 238 4103
rect 204 4001 238 4035
rect 204 3933 238 3967
rect 204 3865 238 3899
rect 204 3797 238 3831
rect 204 3729 238 3763
rect 204 3661 238 3695
rect 646 5565 680 5599
rect 646 5497 680 5531
rect 646 5429 680 5463
rect 646 5361 680 5395
rect 646 5293 680 5327
rect 646 5225 680 5259
rect 646 5157 680 5191
rect 646 5089 680 5123
rect 646 5021 680 5055
rect 646 4953 680 4987
rect 646 4885 680 4919
rect 646 4817 680 4851
rect 646 4749 680 4783
rect 646 4681 680 4715
rect 646 4613 680 4647
rect 646 4545 680 4579
rect 646 4477 680 4511
rect 646 4409 680 4443
rect 646 4341 680 4375
rect 646 4273 680 4307
rect 646 4205 680 4239
rect 646 4137 680 4171
rect 646 4069 680 4103
rect 646 4001 680 4035
rect 646 3933 680 3967
rect 646 3865 680 3899
rect 646 3797 680 3831
rect 646 3729 680 3763
rect 646 3661 680 3695
rect 904 5565 938 5599
rect 904 5497 938 5531
rect 904 5429 938 5463
rect 904 5361 938 5395
rect 904 5293 938 5327
rect 904 5225 938 5259
rect 904 5157 938 5191
rect 904 5089 938 5123
rect 904 5021 938 5055
rect 904 4953 938 4987
rect 904 4885 938 4919
rect 904 4817 938 4851
rect 904 4749 938 4783
rect 904 4681 938 4715
rect 904 4613 938 4647
rect 904 4545 938 4579
rect 904 4477 938 4511
rect 904 4409 938 4443
rect 904 4341 938 4375
rect 904 4273 938 4307
rect 904 4205 938 4239
rect 904 4137 938 4171
rect 904 4069 938 4103
rect 904 4001 938 4035
rect 904 3933 938 3967
rect 904 3865 938 3899
rect 904 3797 938 3831
rect 904 3729 938 3763
rect 904 3661 938 3695
rect 1346 5565 1380 5599
rect 1346 5497 1380 5531
rect 1346 5429 1380 5463
rect 1346 5361 1380 5395
rect 1346 5293 1380 5327
rect 1346 5225 1380 5259
rect 1346 5157 1380 5191
rect 1346 5089 1380 5123
rect 1346 5021 1380 5055
rect 1346 4953 1380 4987
rect 1346 4885 1380 4919
rect 1346 4817 1380 4851
rect 1346 4749 1380 4783
rect 1346 4681 1380 4715
rect 1346 4613 1380 4647
rect 1346 4545 1380 4579
rect 1346 4477 1380 4511
rect 1346 4409 1380 4443
rect 1346 4341 1380 4375
rect 1346 4273 1380 4307
rect 1346 4205 1380 4239
rect 1346 4137 1380 4171
rect 1346 4069 1380 4103
rect 1346 4001 1380 4035
rect 1346 3933 1380 3967
rect 1346 3865 1380 3899
rect 1346 3797 1380 3831
rect 1346 3729 1380 3763
rect 1346 3661 1380 3695
rect 1604 5565 1638 5599
rect 1604 5497 1638 5531
rect 1604 5429 1638 5463
rect 1604 5361 1638 5395
rect 1604 5293 1638 5327
rect 1604 5225 1638 5259
rect 1604 5157 1638 5191
rect 1604 5089 1638 5123
rect 1604 5021 1638 5055
rect 1604 4953 1638 4987
rect 1604 4885 1638 4919
rect 1604 4817 1638 4851
rect 1604 4749 1638 4783
rect 1604 4681 1638 4715
rect 1604 4613 1638 4647
rect 1604 4545 1638 4579
rect 1604 4477 1638 4511
rect 1604 4409 1638 4443
rect 1604 4341 1638 4375
rect 1604 4273 1638 4307
rect 1604 4205 1638 4239
rect 1604 4137 1638 4171
rect 1604 4069 1638 4103
rect 1604 4001 1638 4035
rect 1604 3933 1638 3967
rect 1604 3865 1638 3899
rect 1604 3797 1638 3831
rect 1604 3729 1638 3763
rect 1604 3661 1638 3695
rect 2046 5565 2080 5599
rect 2046 5497 2080 5531
rect 2046 5429 2080 5463
rect 2046 5361 2080 5395
rect 2046 5293 2080 5327
rect 2046 5225 2080 5259
rect 2046 5157 2080 5191
rect 2046 5089 2080 5123
rect 2046 5021 2080 5055
rect 2046 4953 2080 4987
rect 2046 4885 2080 4919
rect 2046 4817 2080 4851
rect 2046 4749 2080 4783
rect 2046 4681 2080 4715
rect 2046 4613 2080 4647
rect 2046 4545 2080 4579
rect 2046 4477 2080 4511
rect 2046 4409 2080 4443
rect 2046 4341 2080 4375
rect 2046 4273 2080 4307
rect 2046 4205 2080 4239
rect 2046 4137 2080 4171
rect 2046 4069 2080 4103
rect 2046 4001 2080 4035
rect 2046 3933 2080 3967
rect 2046 3865 2080 3899
rect 2046 3797 2080 3831
rect 2046 3729 2080 3763
rect 2046 3661 2080 3695
rect 2304 5565 2338 5599
rect 2304 5497 2338 5531
rect 2304 5429 2338 5463
rect 2304 5361 2338 5395
rect 2304 5293 2338 5327
rect 2304 5225 2338 5259
rect 2304 5157 2338 5191
rect 2304 5089 2338 5123
rect 2304 5021 2338 5055
rect 2304 4953 2338 4987
rect 2304 4885 2338 4919
rect 2304 4817 2338 4851
rect 2304 4749 2338 4783
rect 2304 4681 2338 4715
rect 2304 4613 2338 4647
rect 2304 4545 2338 4579
rect 2304 4477 2338 4511
rect 2304 4409 2338 4443
rect 2304 4341 2338 4375
rect 2304 4273 2338 4307
rect 2304 4205 2338 4239
rect 2304 4137 2338 4171
rect 2304 4069 2338 4103
rect 2304 4001 2338 4035
rect 2304 3933 2338 3967
rect 2304 3865 2338 3899
rect 2304 3797 2338 3831
rect 2304 3729 2338 3763
rect 2304 3661 2338 3695
rect 3746 5565 3780 5599
rect 3746 5497 3780 5531
rect 3746 5429 3780 5463
rect 3746 5361 3780 5395
rect 3746 5293 3780 5327
rect 3746 5225 3780 5259
rect 3746 5157 3780 5191
rect 3746 5089 3780 5123
rect 3746 5021 3780 5055
rect 3746 4953 3780 4987
rect 3746 4885 3780 4919
rect 3746 4817 3780 4851
rect 3746 4749 3780 4783
rect 3746 4681 3780 4715
rect 3746 4613 3780 4647
rect 3746 4545 3780 4579
rect 3746 4477 3780 4511
rect 3746 4409 3780 4443
rect 3746 4341 3780 4375
rect 3746 4273 3780 4307
rect 3746 4205 3780 4239
rect 3746 4137 3780 4171
rect 3746 4069 3780 4103
rect 3746 4001 3780 4035
rect 3746 3933 3780 3967
rect 3746 3865 3780 3899
rect 3746 3797 3780 3831
rect 3746 3729 3780 3763
rect 3746 3661 3780 3695
rect 4004 5565 4038 5599
rect 4004 5497 4038 5531
rect 4004 5429 4038 5463
rect 4004 5361 4038 5395
rect 4004 5293 4038 5327
rect 4004 5225 4038 5259
rect 4004 5157 4038 5191
rect 4004 5089 4038 5123
rect 4004 5021 4038 5055
rect 4004 4953 4038 4987
rect 4004 4885 4038 4919
rect 4004 4817 4038 4851
rect 4004 4749 4038 4783
rect 4004 4681 4038 4715
rect 4004 4613 4038 4647
rect 4004 4545 4038 4579
rect 4004 4477 4038 4511
rect 4004 4409 4038 4443
rect 4004 4341 4038 4375
rect 4004 4273 4038 4307
rect 4004 4205 4038 4239
rect 4004 4137 4038 4171
rect 4004 4069 4038 4103
rect 4004 4001 4038 4035
rect 4004 3933 4038 3967
rect 4004 3865 4038 3899
rect 4004 3797 4038 3831
rect 4004 3729 4038 3763
rect 4004 3661 4038 3695
rect 4446 5565 4480 5599
rect 4446 5497 4480 5531
rect 4446 5429 4480 5463
rect 4446 5361 4480 5395
rect 4446 5293 4480 5327
rect 4446 5225 4480 5259
rect 4446 5157 4480 5191
rect 4446 5089 4480 5123
rect 4446 5021 4480 5055
rect 4446 4953 4480 4987
rect 4446 4885 4480 4919
rect 4446 4817 4480 4851
rect 4446 4749 4480 4783
rect 4446 4681 4480 4715
rect 4446 4613 4480 4647
rect 4446 4545 4480 4579
rect 4446 4477 4480 4511
rect 4446 4409 4480 4443
rect 4446 4341 4480 4375
rect 4446 4273 4480 4307
rect 4446 4205 4480 4239
rect 4446 4137 4480 4171
rect 4446 4069 4480 4103
rect 4446 4001 4480 4035
rect 4446 3933 4480 3967
rect 4446 3865 4480 3899
rect 4446 3797 4480 3831
rect 4446 3729 4480 3763
rect 4446 3661 4480 3695
rect 4704 5565 4738 5599
rect 4704 5497 4738 5531
rect 4704 5429 4738 5463
rect 4704 5361 4738 5395
rect 4704 5293 4738 5327
rect 4704 5225 4738 5259
rect 4704 5157 4738 5191
rect 4704 5089 4738 5123
rect 4704 5021 4738 5055
rect 4704 4953 4738 4987
rect 4704 4885 4738 4919
rect 4704 4817 4738 4851
rect 4704 4749 4738 4783
rect 4704 4681 4738 4715
rect 4704 4613 4738 4647
rect 4704 4545 4738 4579
rect 4704 4477 4738 4511
rect 4704 4409 4738 4443
rect 4704 4341 4738 4375
rect 4704 4273 4738 4307
rect 4704 4205 4738 4239
rect 4704 4137 4738 4171
rect 4704 4069 4738 4103
rect 4704 4001 4738 4035
rect 4704 3933 4738 3967
rect 4704 3865 4738 3899
rect 4704 3797 4738 3831
rect 4704 3729 4738 3763
rect 4704 3661 4738 3695
rect 5146 5565 5180 5599
rect 5146 5497 5180 5531
rect 5146 5429 5180 5463
rect 5146 5361 5180 5395
rect 5146 5293 5180 5327
rect 5146 5225 5180 5259
rect 5146 5157 5180 5191
rect 5146 5089 5180 5123
rect 5146 5021 5180 5055
rect 5146 4953 5180 4987
rect 5146 4885 5180 4919
rect 5146 4817 5180 4851
rect 5146 4749 5180 4783
rect 5146 4681 5180 4715
rect 5146 4613 5180 4647
rect 5146 4545 5180 4579
rect 5146 4477 5180 4511
rect 5146 4409 5180 4443
rect 5146 4341 5180 4375
rect 5146 4273 5180 4307
rect 5146 4205 5180 4239
rect 5146 4137 5180 4171
rect 5146 4069 5180 4103
rect 5146 4001 5180 4035
rect 5146 3933 5180 3967
rect 5146 3865 5180 3899
rect 5146 3797 5180 3831
rect 5146 3729 5180 3763
rect 5146 3661 5180 3695
rect 5404 5565 5438 5599
rect 5404 5497 5438 5531
rect 5404 5429 5438 5463
rect 5404 5361 5438 5395
rect 5404 5293 5438 5327
rect 5404 5225 5438 5259
rect 5404 5157 5438 5191
rect 5404 5089 5438 5123
rect 5404 5021 5438 5055
rect 5404 4953 5438 4987
rect 5404 4885 5438 4919
rect 5404 4817 5438 4851
rect 5404 4749 5438 4783
rect 5404 4681 5438 4715
rect 5404 4613 5438 4647
rect 5404 4545 5438 4579
rect 5404 4477 5438 4511
rect 5404 4409 5438 4443
rect 5404 4341 5438 4375
rect 5404 4273 5438 4307
rect 5404 4205 5438 4239
rect 5404 4137 5438 4171
rect 5404 4069 5438 4103
rect 5404 4001 5438 4035
rect 5404 3933 5438 3967
rect 5404 3865 5438 3899
rect 5404 3797 5438 3831
rect 5404 3729 5438 3763
rect 5404 3661 5438 3695
rect 5846 5565 5880 5599
rect 5846 5497 5880 5531
rect 5846 5429 5880 5463
rect 5846 5361 5880 5395
rect 5846 5293 5880 5327
rect 5846 5225 5880 5259
rect 5846 5157 5880 5191
rect 5846 5089 5880 5123
rect 5846 5021 5880 5055
rect 5846 4953 5880 4987
rect 5846 4885 5880 4919
rect 5846 4817 5880 4851
rect 5846 4749 5880 4783
rect 5846 4681 5880 4715
rect 5846 4613 5880 4647
rect 5846 4545 5880 4579
rect 5846 4477 5880 4511
rect 5846 4409 5880 4443
rect 5846 4341 5880 4375
rect 5846 4273 5880 4307
rect 5846 4205 5880 4239
rect 5846 4137 5880 4171
rect 5846 4069 5880 4103
rect 5846 4001 5880 4035
rect 5846 3933 5880 3967
rect 5846 3865 5880 3899
rect 5846 3797 5880 3831
rect 5846 3729 5880 3763
rect 5846 3661 5880 3695
rect 6104 5565 6138 5599
rect 6104 5497 6138 5531
rect 6104 5429 6138 5463
rect 6104 5361 6138 5395
rect 6104 5293 6138 5327
rect 6104 5225 6138 5259
rect 6104 5157 6138 5191
rect 6104 5089 6138 5123
rect 6104 5021 6138 5055
rect 6104 4953 6138 4987
rect 6104 4885 6138 4919
rect 6104 4817 6138 4851
rect 6104 4749 6138 4783
rect 6104 4681 6138 4715
rect 6104 4613 6138 4647
rect 6104 4545 6138 4579
rect 6104 4477 6138 4511
rect 6104 4409 6138 4443
rect 6104 4341 6138 4375
rect 6104 4273 6138 4307
rect 6104 4205 6138 4239
rect 6104 4137 6138 4171
rect 6104 4069 6138 4103
rect 6104 4001 6138 4035
rect 6104 3933 6138 3967
rect 6104 3865 6138 3899
rect 6104 3797 6138 3831
rect 6104 3729 6138 3763
rect 6104 3661 6138 3695
rect 6546 5565 6580 5599
rect 6546 5497 6580 5531
rect 6546 5429 6580 5463
rect 6546 5361 6580 5395
rect 6546 5293 6580 5327
rect 6546 5225 6580 5259
rect 6546 5157 6580 5191
rect 6546 5089 6580 5123
rect 6546 5021 6580 5055
rect 6546 4953 6580 4987
rect 6546 4885 6580 4919
rect 6546 4817 6580 4851
rect 6546 4749 6580 4783
rect 6546 4681 6580 4715
rect 6546 4613 6580 4647
rect 6546 4545 6580 4579
rect 6546 4477 6580 4511
rect 6546 4409 6580 4443
rect 6546 4341 6580 4375
rect 6546 4273 6580 4307
rect 6546 4205 6580 4239
rect 6546 4137 6580 4171
rect 6546 4069 6580 4103
rect 6546 4001 6580 4035
rect 6546 3933 6580 3967
rect 6546 3865 6580 3899
rect 6546 3797 6580 3831
rect 6546 3729 6580 3763
rect 6546 3661 6580 3695
rect 6804 5565 6838 5599
rect 6804 5497 6838 5531
rect 6804 5429 6838 5463
rect 6804 5361 6838 5395
rect 6804 5293 6838 5327
rect 6804 5225 6838 5259
rect 6804 5157 6838 5191
rect 6804 5089 6838 5123
rect 6804 5021 6838 5055
rect 6804 4953 6838 4987
rect 6804 4885 6838 4919
rect 6804 4817 6838 4851
rect 6804 4749 6838 4783
rect 6804 4681 6838 4715
rect 6804 4613 6838 4647
rect 6804 4545 6838 4579
rect 6804 4477 6838 4511
rect 6804 4409 6838 4443
rect 6804 4341 6838 4375
rect 6804 4273 6838 4307
rect 6804 4205 6838 4239
rect 6804 4137 6838 4171
rect 6804 4069 6838 4103
rect 6804 4001 6838 4035
rect 6804 3933 6838 3967
rect 6804 3865 6838 3899
rect 6804 3797 6838 3831
rect 6804 3729 6838 3763
rect 6804 3661 6838 3695
rect 7246 5565 7280 5599
rect 7246 5497 7280 5531
rect 7246 5429 7280 5463
rect 7246 5361 7280 5395
rect 7246 5293 7280 5327
rect 7246 5225 7280 5259
rect 7246 5157 7280 5191
rect 7246 5089 7280 5123
rect 7246 5021 7280 5055
rect 7246 4953 7280 4987
rect 7246 4885 7280 4919
rect 7246 4817 7280 4851
rect 7246 4749 7280 4783
rect 7246 4681 7280 4715
rect 7246 4613 7280 4647
rect 7246 4545 7280 4579
rect 7246 4477 7280 4511
rect 7246 4409 7280 4443
rect 7246 4341 7280 4375
rect 7246 4273 7280 4307
rect 7246 4205 7280 4239
rect 7246 4137 7280 4171
rect 7246 4069 7280 4103
rect 7246 4001 7280 4035
rect 7246 3933 7280 3967
rect 7246 3865 7280 3899
rect 7246 3797 7280 3831
rect 7246 3729 7280 3763
rect 7246 3661 7280 3695
rect 7504 5565 7538 5599
rect 7504 5497 7538 5531
rect 7504 5429 7538 5463
rect 7504 5361 7538 5395
rect 7504 5293 7538 5327
rect 7504 5225 7538 5259
rect 7504 5157 7538 5191
rect 7504 5089 7538 5123
rect 7504 5021 7538 5055
rect 7504 4953 7538 4987
rect 7504 4885 7538 4919
rect 7504 4817 7538 4851
rect 7504 4749 7538 4783
rect 7504 4681 7538 4715
rect 7504 4613 7538 4647
rect 7504 4545 7538 4579
rect 7504 4477 7538 4511
rect 7504 4409 7538 4443
rect 7504 4341 7538 4375
rect 7504 4273 7538 4307
rect 7504 4205 7538 4239
rect 7504 4137 7538 4171
rect 7504 4069 7538 4103
rect 7504 4001 7538 4035
rect 7504 3933 7538 3967
rect 7504 3865 7538 3899
rect 7504 3797 7538 3831
rect 7504 3729 7538 3763
rect 7504 3661 7538 3695
rect 7946 5565 7980 5599
rect 7946 5497 7980 5531
rect 7946 5429 7980 5463
rect 7946 5361 7980 5395
rect 7946 5293 7980 5327
rect 7946 5225 7980 5259
rect 7946 5157 7980 5191
rect 7946 5089 7980 5123
rect 7946 5021 7980 5055
rect 7946 4953 7980 4987
rect 7946 4885 7980 4919
rect 7946 4817 7980 4851
rect 7946 4749 7980 4783
rect 7946 4681 7980 4715
rect 7946 4613 7980 4647
rect 7946 4545 7980 4579
rect 7946 4477 7980 4511
rect 7946 4409 7980 4443
rect 7946 4341 7980 4375
rect 7946 4273 7980 4307
rect 7946 4205 7980 4239
rect 7946 4137 7980 4171
rect 7946 4069 7980 4103
rect 7946 4001 7980 4035
rect 7946 3933 7980 3967
rect 7946 3865 7980 3899
rect 7946 3797 7980 3831
rect 7946 3729 7980 3763
rect 7946 3661 7980 3695
rect 8204 5565 8238 5599
rect 8204 5497 8238 5531
rect 8204 5429 8238 5463
rect 8204 5361 8238 5395
rect 8204 5293 8238 5327
rect 8204 5225 8238 5259
rect 8204 5157 8238 5191
rect 8204 5089 8238 5123
rect 8204 5021 8238 5055
rect 8204 4953 8238 4987
rect 8204 4885 8238 4919
rect 8204 4817 8238 4851
rect 8204 4749 8238 4783
rect 8204 4681 8238 4715
rect 8204 4613 8238 4647
rect 8204 4545 8238 4579
rect 8204 4477 8238 4511
rect 8204 4409 8238 4443
rect 8204 4341 8238 4375
rect 8204 4273 8238 4307
rect 8204 4205 8238 4239
rect 8204 4137 8238 4171
rect 8204 4069 8238 4103
rect 8204 4001 8238 4035
rect 8204 3933 8238 3967
rect 8204 3865 8238 3899
rect 8204 3797 8238 3831
rect 8204 3729 8238 3763
rect 8204 3661 8238 3695
rect 8646 5565 8680 5599
rect 8646 5497 8680 5531
rect 8646 5429 8680 5463
rect 8646 5361 8680 5395
rect 8646 5293 8680 5327
rect 8646 5225 8680 5259
rect 8646 5157 8680 5191
rect 8646 5089 8680 5123
rect 8646 5021 8680 5055
rect 8646 4953 8680 4987
rect 8646 4885 8680 4919
rect 8646 4817 8680 4851
rect 8646 4749 8680 4783
rect 8646 4681 8680 4715
rect 8646 4613 8680 4647
rect 8646 4545 8680 4579
rect 8646 4477 8680 4511
rect 8646 4409 8680 4443
rect 8646 4341 8680 4375
rect 8646 4273 8680 4307
rect 8646 4205 8680 4239
rect 8646 4137 8680 4171
rect 8646 4069 8680 4103
rect 8646 4001 8680 4035
rect 8646 3933 8680 3967
rect 8646 3865 8680 3899
rect 8646 3797 8680 3831
rect 8646 3729 8680 3763
rect 8646 3661 8680 3695
rect 8904 5565 8938 5599
rect 8904 5497 8938 5531
rect 8904 5429 8938 5463
rect 8904 5361 8938 5395
rect 8904 5293 8938 5327
rect 8904 5225 8938 5259
rect 8904 5157 8938 5191
rect 8904 5089 8938 5123
rect 8904 5021 8938 5055
rect 8904 4953 8938 4987
rect 8904 4885 8938 4919
rect 8904 4817 8938 4851
rect 8904 4749 8938 4783
rect 8904 4681 8938 4715
rect 8904 4613 8938 4647
rect 8904 4545 8938 4579
rect 8904 4477 8938 4511
rect 8904 4409 8938 4443
rect 8904 4341 8938 4375
rect 8904 4273 8938 4307
rect 8904 4205 8938 4239
rect 8904 4137 8938 4171
rect 8904 4069 8938 4103
rect 8904 4001 8938 4035
rect 8904 3933 8938 3967
rect 8904 3865 8938 3899
rect 8904 3797 8938 3831
rect 8904 3729 8938 3763
rect 8904 3661 8938 3695
rect 9346 5565 9380 5599
rect 9346 5497 9380 5531
rect 9346 5429 9380 5463
rect 9346 5361 9380 5395
rect 9346 5293 9380 5327
rect 9346 5225 9380 5259
rect 9346 5157 9380 5191
rect 9346 5089 9380 5123
rect 9346 5021 9380 5055
rect 9346 4953 9380 4987
rect 9346 4885 9380 4919
rect 9346 4817 9380 4851
rect 9346 4749 9380 4783
rect 9346 4681 9380 4715
rect 9346 4613 9380 4647
rect 9346 4545 9380 4579
rect 9346 4477 9380 4511
rect 9346 4409 9380 4443
rect 9346 4341 9380 4375
rect 9346 4273 9380 4307
rect 9346 4205 9380 4239
rect 9346 4137 9380 4171
rect 9346 4069 9380 4103
rect 9346 4001 9380 4035
rect 9346 3933 9380 3967
rect 9346 3865 9380 3899
rect 9346 3797 9380 3831
rect 9346 3729 9380 3763
rect 9346 3661 9380 3695
rect 9604 5565 9638 5599
rect 9604 5497 9638 5531
rect 9604 5429 9638 5463
rect 9604 5361 9638 5395
rect 9604 5293 9638 5327
rect 9604 5225 9638 5259
rect 9604 5157 9638 5191
rect 9604 5089 9638 5123
rect 9604 5021 9638 5055
rect 9604 4953 9638 4987
rect 9604 4885 9638 4919
rect 9604 4817 9638 4851
rect 9604 4749 9638 4783
rect 9604 4681 9638 4715
rect 9604 4613 9638 4647
rect 9604 4545 9638 4579
rect 9604 4477 9638 4511
rect 9604 4409 9638 4443
rect 9604 4341 9638 4375
rect 9604 4273 9638 4307
rect 9604 4205 9638 4239
rect 9604 4137 9638 4171
rect 9604 4069 9638 4103
rect 9604 4001 9638 4035
rect 9604 3933 9638 3967
rect 9604 3865 9638 3899
rect 9604 3797 9638 3831
rect 9604 3729 9638 3763
rect 9604 3661 9638 3695
rect 10046 5565 10080 5599
rect 10046 5497 10080 5531
rect 10046 5429 10080 5463
rect 10046 5361 10080 5395
rect 10046 5293 10080 5327
rect 10046 5225 10080 5259
rect 10046 5157 10080 5191
rect 10046 5089 10080 5123
rect 10046 5021 10080 5055
rect 10046 4953 10080 4987
rect 10046 4885 10080 4919
rect 10046 4817 10080 4851
rect 10046 4749 10080 4783
rect 10046 4681 10080 4715
rect 10046 4613 10080 4647
rect 10046 4545 10080 4579
rect 10046 4477 10080 4511
rect 10046 4409 10080 4443
rect 10046 4341 10080 4375
rect 10046 4273 10080 4307
rect 10046 4205 10080 4239
rect 10046 4137 10080 4171
rect 10046 4069 10080 4103
rect 10046 4001 10080 4035
rect 10046 3933 10080 3967
rect 10046 3865 10080 3899
rect 10046 3797 10080 3831
rect 10046 3729 10080 3763
rect 10046 3661 10080 3695
rect 10304 5565 10338 5599
rect 10304 5497 10338 5531
rect 10304 5429 10338 5463
rect 10304 5361 10338 5395
rect 10304 5293 10338 5327
rect 10304 5225 10338 5259
rect 10304 5157 10338 5191
rect 10304 5089 10338 5123
rect 10304 5021 10338 5055
rect 10304 4953 10338 4987
rect 10304 4885 10338 4919
rect 10304 4817 10338 4851
rect 10304 4749 10338 4783
rect 10304 4681 10338 4715
rect 10304 4613 10338 4647
rect 10304 4545 10338 4579
rect 10304 4477 10338 4511
rect 10304 4409 10338 4443
rect 10304 4341 10338 4375
rect 10304 4273 10338 4307
rect 10304 4205 10338 4239
rect 10304 4137 10338 4171
rect 10304 4069 10338 4103
rect 10304 4001 10338 4035
rect 10304 3933 10338 3967
rect 10304 3865 10338 3899
rect 10304 3797 10338 3831
rect 10304 3729 10338 3763
rect 10304 3661 10338 3695
rect 1088 1867 1122 1901
rect 1088 1799 1122 1833
rect 1088 1731 1122 1765
rect 1546 1867 1580 1901
rect 1546 1799 1580 1833
rect 1546 1731 1580 1765
rect 2088 1867 2122 1901
rect 2088 1799 2122 1833
rect 2088 1731 2122 1765
rect 2546 1867 2580 1901
rect 2546 1799 2580 1833
rect 2546 1731 2580 1765
rect 3088 1867 3122 1901
rect 3088 1799 3122 1833
rect 3088 1731 3122 1765
rect 3546 1867 3580 1901
rect 3546 1799 3580 1833
rect 3546 1731 3580 1765
rect 4088 1867 4122 1901
rect 4088 1799 4122 1833
rect 4088 1731 4122 1765
rect 4546 1867 4580 1901
rect 4546 1799 4580 1833
rect 4546 1731 4580 1765
rect 5088 1867 5122 1901
rect 5088 1799 5122 1833
rect 5088 1731 5122 1765
rect 5546 1867 5580 1901
rect 5546 1799 5580 1833
rect 5546 1731 5580 1765
rect 6088 1867 6122 1901
rect 6088 1799 6122 1833
rect 6088 1731 6122 1765
rect 6546 1867 6580 1901
rect 6546 1799 6580 1833
rect 6546 1731 6580 1765
rect 7088 1867 7122 1901
rect 7088 1799 7122 1833
rect 7088 1731 7122 1765
rect 7546 1867 7580 1901
rect 7546 1799 7580 1833
rect 7546 1731 7580 1765
rect 8088 1867 8122 1901
rect 8088 1799 8122 1833
rect 8088 1731 8122 1765
rect 8546 1867 8580 1901
rect 8546 1799 8580 1833
rect 8546 1731 8580 1765
rect 9088 1867 9122 1901
rect 9088 1799 9122 1833
rect 9088 1731 9122 1765
rect 9546 1867 9580 1901
rect 9546 1799 9580 1833
rect 9546 1731 9580 1765
rect 10088 1867 10122 1901
rect 10088 1799 10122 1833
rect 10088 1731 10122 1765
rect 10546 1867 10580 1901
rect 10546 1799 10580 1833
rect 10546 1731 10580 1765
rect 1088 1367 1122 1401
rect 1088 1299 1122 1333
rect 1088 1231 1122 1265
rect 1546 1367 1580 1401
rect 1546 1299 1580 1333
rect 1546 1231 1580 1265
rect 2088 1367 2122 1401
rect 2088 1299 2122 1333
rect 2088 1231 2122 1265
rect 2546 1367 2580 1401
rect 2546 1299 2580 1333
rect 2546 1231 2580 1265
rect 3088 1367 3122 1401
rect 3088 1299 3122 1333
rect 3088 1231 3122 1265
rect 3546 1367 3580 1401
rect 3546 1299 3580 1333
rect 3546 1231 3580 1265
rect 4088 1367 4122 1401
rect 4088 1299 4122 1333
rect 4088 1231 4122 1265
rect 4546 1367 4580 1401
rect 4546 1299 4580 1333
rect 4546 1231 4580 1265
rect 5088 1367 5122 1401
rect 5088 1299 5122 1333
rect 5088 1231 5122 1265
rect 5546 1367 5580 1401
rect 5546 1299 5580 1333
rect 5546 1231 5580 1265
rect 6088 1367 6122 1401
rect 6088 1299 6122 1333
rect 6088 1231 6122 1265
rect 6546 1367 6580 1401
rect 6546 1299 6580 1333
rect 6546 1231 6580 1265
rect 7088 1367 7122 1401
rect 7088 1299 7122 1333
rect 7088 1231 7122 1265
rect 7546 1367 7580 1401
rect 7546 1299 7580 1333
rect 7546 1231 7580 1265
rect 8088 1367 8122 1401
rect 8088 1299 8122 1333
rect 8088 1231 8122 1265
rect 8546 1367 8580 1401
rect 8546 1299 8580 1333
rect 8546 1231 8580 1265
rect 9088 1367 9122 1401
rect 9088 1299 9122 1333
rect 9088 1231 9122 1265
rect 9546 1367 9580 1401
rect 9546 1299 9580 1333
rect 9546 1231 9580 1265
rect 10088 1367 10122 1401
rect 10088 1299 10122 1333
rect 10088 1231 10122 1265
rect 10546 1367 10580 1401
rect 10546 1299 10580 1333
rect 10546 1231 10580 1265
<< mvpdiffc >>
rect 1978 8462 2012 8496
rect 1978 8394 2012 8428
rect 1978 8326 2012 8360
rect 1978 8258 2012 8292
rect 1978 8190 2012 8224
rect 1978 8122 2012 8156
rect 2436 8462 2470 8496
rect 2436 8394 2470 8428
rect 2436 8326 2470 8360
rect 2436 8258 2470 8292
rect 2436 8190 2470 8224
rect 2436 8122 2470 8156
rect 2978 8462 3012 8496
rect 2978 8394 3012 8428
rect 2978 8326 3012 8360
rect 2978 8258 3012 8292
rect 2978 8190 3012 8224
rect 2978 8122 3012 8156
rect 3436 8462 3470 8496
rect 3436 8394 3470 8428
rect 3436 8326 3470 8360
rect 3436 8258 3470 8292
rect 3436 8190 3470 8224
rect 3436 8122 3470 8156
rect 1978 7722 2012 7756
rect 1978 7654 2012 7688
rect 1978 7586 2012 7620
rect 1978 7518 2012 7552
rect 1978 7450 2012 7484
rect 1978 7382 2012 7416
rect 2436 7722 2470 7756
rect 2436 7654 2470 7688
rect 2436 7586 2470 7620
rect 2436 7518 2470 7552
rect 2436 7450 2470 7484
rect 2436 7382 2470 7416
rect 2978 7722 3012 7756
rect 2978 7654 3012 7688
rect 2978 7586 3012 7620
rect 2978 7518 3012 7552
rect 2978 7450 3012 7484
rect 2978 7382 3012 7416
rect 3436 7722 3470 7756
rect 3436 7654 3470 7688
rect 3436 7586 3470 7620
rect 3436 7518 3470 7552
rect 3436 7450 3470 7484
rect 3436 7382 3470 7416
rect 11696 6802 11730 6836
rect 11696 6734 11730 6768
rect 11696 6666 11730 6700
rect 11696 6598 11730 6632
rect 11696 6530 11730 6564
rect 11696 6462 11730 6496
rect 12154 6802 12188 6836
rect 12154 6734 12188 6768
rect 12154 6666 12188 6700
rect 12154 6598 12188 6632
rect 12154 6530 12188 6564
rect 12154 6462 12188 6496
rect 12596 6802 12630 6836
rect 12596 6734 12630 6768
rect 12596 6666 12630 6700
rect 12596 6598 12630 6632
rect 12596 6530 12630 6564
rect 12596 6462 12630 6496
rect 13054 6802 13088 6836
rect 13054 6734 13088 6768
rect 13054 6666 13088 6700
rect 13054 6598 13088 6632
rect 13054 6530 13088 6564
rect 13054 6462 13088 6496
rect 13496 6802 13530 6836
rect 13496 6734 13530 6768
rect 13496 6666 13530 6700
rect 13496 6598 13530 6632
rect 13496 6530 13530 6564
rect 13496 6462 13530 6496
rect 13954 6802 13988 6836
rect 13954 6734 13988 6768
rect 13954 6666 13988 6700
rect 13954 6598 13988 6632
rect 13954 6530 13988 6564
rect 13954 6462 13988 6496
rect 14396 6802 14430 6836
rect 14396 6734 14430 6768
rect 14396 6666 14430 6700
rect 14396 6598 14430 6632
rect 14396 6530 14430 6564
rect 14396 6462 14430 6496
rect 14854 6802 14888 6836
rect 14854 6734 14888 6768
rect 14854 6666 14888 6700
rect 14854 6598 14888 6632
rect 14854 6530 14888 6564
rect 14854 6462 14888 6496
rect 15296 6802 15330 6836
rect 15296 6734 15330 6768
rect 15296 6666 15330 6700
rect 15296 6598 15330 6632
rect 15296 6530 15330 6564
rect 15296 6462 15330 6496
rect 15754 6802 15788 6836
rect 15754 6734 15788 6768
rect 15754 6666 15788 6700
rect 15754 6598 15788 6632
rect 15754 6530 15788 6564
rect 15754 6462 15788 6496
rect 16196 6802 16230 6836
rect 16196 6734 16230 6768
rect 16196 6666 16230 6700
rect 16196 6598 16230 6632
rect 16196 6530 16230 6564
rect 16196 6462 16230 6496
rect 16654 6802 16688 6836
rect 16654 6734 16688 6768
rect 16654 6666 16688 6700
rect 16654 6598 16688 6632
rect 16654 6530 16688 6564
rect 16654 6462 16688 6496
rect 17096 6802 17130 6836
rect 17096 6734 17130 6768
rect 17096 6666 17130 6700
rect 17096 6598 17130 6632
rect 17096 6530 17130 6564
rect 17096 6462 17130 6496
rect 17554 6802 17588 6836
rect 17554 6734 17588 6768
rect 17554 6666 17588 6700
rect 17554 6598 17588 6632
rect 17554 6530 17588 6564
rect 17554 6462 17588 6496
rect 17996 6802 18030 6836
rect 17996 6734 18030 6768
rect 17996 6666 18030 6700
rect 17996 6598 18030 6632
rect 17996 6530 18030 6564
rect 17996 6462 18030 6496
rect 18454 6802 18488 6836
rect 18454 6734 18488 6768
rect 18454 6666 18488 6700
rect 18454 6598 18488 6632
rect 18454 6530 18488 6564
rect 18454 6462 18488 6496
rect 11696 6062 11730 6096
rect 11696 5994 11730 6028
rect 11696 5926 11730 5960
rect 11696 5858 11730 5892
rect 11696 5790 11730 5824
rect 11696 5722 11730 5756
rect 12154 6062 12188 6096
rect 12154 5994 12188 6028
rect 12154 5926 12188 5960
rect 12154 5858 12188 5892
rect 12154 5790 12188 5824
rect 12154 5722 12188 5756
rect 12596 6062 12630 6096
rect 12596 5994 12630 6028
rect 12596 5926 12630 5960
rect 12596 5858 12630 5892
rect 12596 5790 12630 5824
rect 12596 5722 12630 5756
rect 13054 6062 13088 6096
rect 13054 5994 13088 6028
rect 13054 5926 13088 5960
rect 13054 5858 13088 5892
rect 13054 5790 13088 5824
rect 13054 5722 13088 5756
rect 13496 6062 13530 6096
rect 13496 5994 13530 6028
rect 13496 5926 13530 5960
rect 13496 5858 13530 5892
rect 13496 5790 13530 5824
rect 13496 5722 13530 5756
rect 13954 6062 13988 6096
rect 13954 5994 13988 6028
rect 13954 5926 13988 5960
rect 13954 5858 13988 5892
rect 13954 5790 13988 5824
rect 13954 5722 13988 5756
rect 14396 6062 14430 6096
rect 14396 5994 14430 6028
rect 14396 5926 14430 5960
rect 14396 5858 14430 5892
rect 14396 5790 14430 5824
rect 14396 5722 14430 5756
rect 14854 6062 14888 6096
rect 14854 5994 14888 6028
rect 14854 5926 14888 5960
rect 14854 5858 14888 5892
rect 14854 5790 14888 5824
rect 14854 5722 14888 5756
rect 15296 6062 15330 6096
rect 15296 5994 15330 6028
rect 15296 5926 15330 5960
rect 15296 5858 15330 5892
rect 15296 5790 15330 5824
rect 15296 5722 15330 5756
rect 15754 6062 15788 6096
rect 15754 5994 15788 6028
rect 15754 5926 15788 5960
rect 15754 5858 15788 5892
rect 15754 5790 15788 5824
rect 15754 5722 15788 5756
rect 16196 6062 16230 6096
rect 16196 5994 16230 6028
rect 16196 5926 16230 5960
rect 16196 5858 16230 5892
rect 16196 5790 16230 5824
rect 16196 5722 16230 5756
rect 16654 6062 16688 6096
rect 16654 5994 16688 6028
rect 16654 5926 16688 5960
rect 16654 5858 16688 5892
rect 16654 5790 16688 5824
rect 16654 5722 16688 5756
rect 17096 6062 17130 6096
rect 17096 5994 17130 6028
rect 17096 5926 17130 5960
rect 17096 5858 17130 5892
rect 17096 5790 17130 5824
rect 17096 5722 17130 5756
rect 17554 6062 17588 6096
rect 17554 5994 17588 6028
rect 17554 5926 17588 5960
rect 17554 5858 17588 5892
rect 17554 5790 17588 5824
rect 17554 5722 17588 5756
rect 17996 6062 18030 6096
rect 17996 5994 18030 6028
rect 17996 5926 18030 5960
rect 17996 5858 18030 5892
rect 17996 5790 18030 5824
rect 17996 5722 18030 5756
rect 18454 6062 18488 6096
rect 18454 5994 18488 6028
rect 18454 5926 18488 5960
rect 18454 5858 18488 5892
rect 18454 5790 18488 5824
rect 18454 5722 18488 5756
<< psubdiff >>
rect 21073 7603 21155 7627
rect 21073 7569 21097 7603
rect 21131 7569 21155 7603
rect 21073 7531 21155 7569
rect 21073 7497 21097 7531
rect 21131 7497 21155 7531
rect 21073 7473 21155 7497
rect -4176 5925 -4022 5949
rect -4176 5891 -4152 5925
rect -4118 5891 -4080 5925
rect -4046 5891 -4022 5925
rect -4176 5867 -4022 5891
rect -3476 5925 -3322 5949
rect -3476 5891 -3452 5925
rect -3418 5891 -3380 5925
rect -3346 5891 -3322 5925
rect -3476 5867 -3322 5891
rect -2776 5925 -2622 5949
rect -2776 5891 -2752 5925
rect -2718 5891 -2680 5925
rect -2646 5891 -2622 5925
rect -2776 5867 -2622 5891
rect -2076 5925 -1922 5949
rect -2076 5891 -2052 5925
rect -2018 5891 -1980 5925
rect -1946 5891 -1922 5925
rect -2076 5867 -1922 5891
rect -1376 5925 -1222 5949
rect -1376 5891 -1352 5925
rect -1318 5891 -1280 5925
rect -1246 5891 -1222 5925
rect -1376 5867 -1222 5891
rect -676 5925 -522 5949
rect -676 5891 -652 5925
rect -618 5891 -580 5925
rect -546 5891 -522 5925
rect -676 5867 -522 5891
rect 24 5925 178 5949
rect 24 5891 48 5925
rect 82 5891 120 5925
rect 154 5891 178 5925
rect 24 5867 178 5891
rect 724 5925 878 5949
rect 724 5891 748 5925
rect 782 5891 820 5925
rect 854 5891 878 5925
rect 724 5867 878 5891
rect 1424 5925 1578 5949
rect 1424 5891 1448 5925
rect 1482 5891 1520 5925
rect 1554 5891 1578 5925
rect 1424 5867 1578 5891
rect 2124 5925 2278 5949
rect 2124 5891 2148 5925
rect 2182 5891 2220 5925
rect 2254 5891 2278 5925
rect 2124 5867 2278 5891
rect 3824 5925 3978 5949
rect 3824 5891 3848 5925
rect 3882 5891 3920 5925
rect 3954 5891 3978 5925
rect 3824 5867 3978 5891
rect 4524 5925 4678 5949
rect 4524 5891 4548 5925
rect 4582 5891 4620 5925
rect 4654 5891 4678 5925
rect 4524 5867 4678 5891
rect 5224 5925 5378 5949
rect 5224 5891 5248 5925
rect 5282 5891 5320 5925
rect 5354 5891 5378 5925
rect 5224 5867 5378 5891
rect 5924 5925 6078 5949
rect 5924 5891 5948 5925
rect 5982 5891 6020 5925
rect 6054 5891 6078 5925
rect 5924 5867 6078 5891
rect 6624 5925 6778 5949
rect 6624 5891 6648 5925
rect 6682 5891 6720 5925
rect 6754 5891 6778 5925
rect 6624 5867 6778 5891
rect 7324 5925 7478 5949
rect 7324 5891 7348 5925
rect 7382 5891 7420 5925
rect 7454 5891 7478 5925
rect 7324 5867 7478 5891
rect 8024 5925 8178 5949
rect 8024 5891 8048 5925
rect 8082 5891 8120 5925
rect 8154 5891 8178 5925
rect 8024 5867 8178 5891
rect 8724 5925 8878 5949
rect 8724 5891 8748 5925
rect 8782 5891 8820 5925
rect 8854 5891 8878 5925
rect 8724 5867 8878 5891
rect 9424 5925 9578 5949
rect 9424 5891 9448 5925
rect 9482 5891 9520 5925
rect 9554 5891 9578 5925
rect 9424 5867 9578 5891
rect 10124 5925 10278 5949
rect 10124 5891 10148 5925
rect 10182 5891 10220 5925
rect 10254 5891 10278 5925
rect 10124 5867 10278 5891
rect 1261 2134 1415 2158
rect 1261 2100 1285 2134
rect 1319 2100 1357 2134
rect 1391 2100 1415 2134
rect 1261 2076 1415 2100
rect 2261 2134 2415 2158
rect 2261 2100 2285 2134
rect 2319 2100 2357 2134
rect 2391 2100 2415 2134
rect 2261 2076 2415 2100
rect 3261 2134 3415 2158
rect 3261 2100 3285 2134
rect 3319 2100 3357 2134
rect 3391 2100 3415 2134
rect 3261 2076 3415 2100
rect 4261 2134 4415 2158
rect 4261 2100 4285 2134
rect 4319 2100 4357 2134
rect 4391 2100 4415 2134
rect 4261 2076 4415 2100
rect 5261 2134 5415 2158
rect 5261 2100 5285 2134
rect 5319 2100 5357 2134
rect 5391 2100 5415 2134
rect 5261 2076 5415 2100
rect 6261 2134 6415 2158
rect 6261 2100 6285 2134
rect 6319 2100 6357 2134
rect 6391 2100 6415 2134
rect 6261 2076 6415 2100
rect 7261 2134 7415 2158
rect 7261 2100 7285 2134
rect 7319 2100 7357 2134
rect 7391 2100 7415 2134
rect 7261 2076 7415 2100
rect 8261 2134 8415 2158
rect 8261 2100 8285 2134
rect 8319 2100 8357 2134
rect 8391 2100 8415 2134
rect 8261 2076 8415 2100
rect 9261 2134 9415 2158
rect 9261 2100 9285 2134
rect 9319 2100 9357 2134
rect 9391 2100 9415 2134
rect 9261 2076 9415 2100
rect 10261 2134 10415 2158
rect 10261 2100 10285 2134
rect 10319 2100 10357 2134
rect 10391 2100 10415 2134
rect 10261 2076 10415 2100
rect 1260 997 1414 1021
rect 1260 963 1284 997
rect 1318 963 1356 997
rect 1390 963 1414 997
rect 1260 939 1414 963
rect 2260 997 2414 1021
rect 2260 963 2284 997
rect 2318 963 2356 997
rect 2390 963 2414 997
rect 2260 939 2414 963
rect 3260 997 3414 1021
rect 3260 963 3284 997
rect 3318 963 3356 997
rect 3390 963 3414 997
rect 3260 939 3414 963
rect 4260 997 4414 1021
rect 4260 963 4284 997
rect 4318 963 4356 997
rect 4390 963 4414 997
rect 4260 939 4414 963
rect 5260 997 5414 1021
rect 5260 963 5284 997
rect 5318 963 5356 997
rect 5390 963 5414 997
rect 5260 939 5414 963
rect 6260 997 6414 1021
rect 6260 963 6284 997
rect 6318 963 6356 997
rect 6390 963 6414 997
rect 6260 939 6414 963
rect 7260 997 7414 1021
rect 7260 963 7284 997
rect 7318 963 7356 997
rect 7390 963 7414 997
rect 7260 939 7414 963
rect 8260 997 8414 1021
rect 8260 963 8284 997
rect 8318 963 8356 997
rect 8390 963 8414 997
rect 8260 939 8414 963
rect 9260 997 9414 1021
rect 9260 963 9284 997
rect 9318 963 9356 997
rect 9390 963 9414 997
rect 9260 939 9414 963
rect 10260 997 10414 1021
rect 10260 963 10284 997
rect 10318 963 10356 997
rect 10390 963 10414 997
rect 10260 939 10414 963
<< nsubdiff >>
rect 2143 8754 2297 8778
rect 2143 8720 2167 8754
rect 2201 8720 2239 8754
rect 2273 8720 2297 8754
rect 2143 8696 2297 8720
rect 3143 8754 3297 8778
rect 3143 8720 3167 8754
rect 3201 8720 3239 8754
rect 3273 8720 3297 8754
rect 3143 8696 3297 8720
rect 2140 7149 2294 7173
rect 2140 7115 2164 7149
rect 2198 7115 2236 7149
rect 2270 7115 2294 7149
rect 2140 7091 2294 7115
rect 3140 7149 3294 7173
rect 3140 7115 3164 7149
rect 3198 7115 3236 7149
rect 3270 7115 3294 7149
rect 3140 7091 3294 7115
rect 11861 7094 12015 7118
rect 11861 7060 11885 7094
rect 11919 7060 11957 7094
rect 11991 7060 12015 7094
rect 11861 7036 12015 7060
rect 12761 7094 12915 7118
rect 12761 7060 12785 7094
rect 12819 7060 12857 7094
rect 12891 7060 12915 7094
rect 12761 7036 12915 7060
rect 13661 7094 13815 7118
rect 13661 7060 13685 7094
rect 13719 7060 13757 7094
rect 13791 7060 13815 7094
rect 13661 7036 13815 7060
rect 14561 7094 14715 7118
rect 14561 7060 14585 7094
rect 14619 7060 14657 7094
rect 14691 7060 14715 7094
rect 14561 7036 14715 7060
rect 15461 7094 15615 7118
rect 15461 7060 15485 7094
rect 15519 7060 15557 7094
rect 15591 7060 15615 7094
rect 15461 7036 15615 7060
rect 16361 7094 16515 7118
rect 16361 7060 16385 7094
rect 16419 7060 16457 7094
rect 16491 7060 16515 7094
rect 16361 7036 16515 7060
rect 17261 7094 17415 7118
rect 17261 7060 17285 7094
rect 17319 7060 17357 7094
rect 17391 7060 17415 7094
rect 17261 7036 17415 7060
rect 18161 7094 18315 7118
rect 18161 7060 18185 7094
rect 18219 7060 18257 7094
rect 18291 7060 18315 7094
rect 18161 7036 18315 7060
rect 11858 5489 12012 5513
rect 11858 5455 11882 5489
rect 11916 5455 11954 5489
rect 11988 5455 12012 5489
rect 11858 5431 12012 5455
rect 12758 5489 12912 5513
rect 12758 5455 12782 5489
rect 12816 5455 12854 5489
rect 12888 5455 12912 5489
rect 12758 5431 12912 5455
rect 13658 5489 13812 5513
rect 13658 5455 13682 5489
rect 13716 5455 13754 5489
rect 13788 5455 13812 5489
rect 13658 5431 13812 5455
rect 14558 5489 14712 5513
rect 14558 5455 14582 5489
rect 14616 5455 14654 5489
rect 14688 5455 14712 5489
rect 14558 5431 14712 5455
rect 15458 5489 15612 5513
rect 15458 5455 15482 5489
rect 15516 5455 15554 5489
rect 15588 5455 15612 5489
rect 15458 5431 15612 5455
rect 16358 5489 16512 5513
rect 16358 5455 16382 5489
rect 16416 5455 16454 5489
rect 16488 5455 16512 5489
rect 16358 5431 16512 5455
rect 17258 5489 17412 5513
rect 17258 5455 17282 5489
rect 17316 5455 17354 5489
rect 17388 5455 17412 5489
rect 17258 5431 17412 5455
rect 18158 5489 18312 5513
rect 18158 5455 18182 5489
rect 18216 5455 18254 5489
rect 18288 5455 18312 5489
rect 18158 5431 18312 5455
<< psubdiffcont >>
rect 21097 7569 21131 7603
rect 21097 7497 21131 7531
rect -4152 5891 -4118 5925
rect -4080 5891 -4046 5925
rect -3452 5891 -3418 5925
rect -3380 5891 -3346 5925
rect -2752 5891 -2718 5925
rect -2680 5891 -2646 5925
rect -2052 5891 -2018 5925
rect -1980 5891 -1946 5925
rect -1352 5891 -1318 5925
rect -1280 5891 -1246 5925
rect -652 5891 -618 5925
rect -580 5891 -546 5925
rect 48 5891 82 5925
rect 120 5891 154 5925
rect 748 5891 782 5925
rect 820 5891 854 5925
rect 1448 5891 1482 5925
rect 1520 5891 1554 5925
rect 2148 5891 2182 5925
rect 2220 5891 2254 5925
rect 3848 5891 3882 5925
rect 3920 5891 3954 5925
rect 4548 5891 4582 5925
rect 4620 5891 4654 5925
rect 5248 5891 5282 5925
rect 5320 5891 5354 5925
rect 5948 5891 5982 5925
rect 6020 5891 6054 5925
rect 6648 5891 6682 5925
rect 6720 5891 6754 5925
rect 7348 5891 7382 5925
rect 7420 5891 7454 5925
rect 8048 5891 8082 5925
rect 8120 5891 8154 5925
rect 8748 5891 8782 5925
rect 8820 5891 8854 5925
rect 9448 5891 9482 5925
rect 9520 5891 9554 5925
rect 10148 5891 10182 5925
rect 10220 5891 10254 5925
rect 1285 2100 1319 2134
rect 1357 2100 1391 2134
rect 2285 2100 2319 2134
rect 2357 2100 2391 2134
rect 3285 2100 3319 2134
rect 3357 2100 3391 2134
rect 4285 2100 4319 2134
rect 4357 2100 4391 2134
rect 5285 2100 5319 2134
rect 5357 2100 5391 2134
rect 6285 2100 6319 2134
rect 6357 2100 6391 2134
rect 7285 2100 7319 2134
rect 7357 2100 7391 2134
rect 8285 2100 8319 2134
rect 8357 2100 8391 2134
rect 9285 2100 9319 2134
rect 9357 2100 9391 2134
rect 10285 2100 10319 2134
rect 10357 2100 10391 2134
rect 1284 963 1318 997
rect 1356 963 1390 997
rect 2284 963 2318 997
rect 2356 963 2390 997
rect 3284 963 3318 997
rect 3356 963 3390 997
rect 4284 963 4318 997
rect 4356 963 4390 997
rect 5284 963 5318 997
rect 5356 963 5390 997
rect 6284 963 6318 997
rect 6356 963 6390 997
rect 7284 963 7318 997
rect 7356 963 7390 997
rect 8284 963 8318 997
rect 8356 963 8390 997
rect 9284 963 9318 997
rect 9356 963 9390 997
rect 10284 963 10318 997
rect 10356 963 10390 997
<< nsubdiffcont >>
rect 2167 8720 2201 8754
rect 2239 8720 2273 8754
rect 3167 8720 3201 8754
rect 3239 8720 3273 8754
rect 2164 7115 2198 7149
rect 2236 7115 2270 7149
rect 3164 7115 3198 7149
rect 3236 7115 3270 7149
rect 11885 7060 11919 7094
rect 11957 7060 11991 7094
rect 12785 7060 12819 7094
rect 12857 7060 12891 7094
rect 13685 7060 13719 7094
rect 13757 7060 13791 7094
rect 14585 7060 14619 7094
rect 14657 7060 14691 7094
rect 15485 7060 15519 7094
rect 15557 7060 15591 7094
rect 16385 7060 16419 7094
rect 16457 7060 16491 7094
rect 17285 7060 17319 7094
rect 17357 7060 17391 7094
rect 18185 7060 18219 7094
rect 18257 7060 18291 7094
rect 11882 5455 11916 5489
rect 11954 5455 11988 5489
rect 12782 5455 12816 5489
rect 12854 5455 12888 5489
rect 13682 5455 13716 5489
rect 13754 5455 13788 5489
rect 14582 5455 14616 5489
rect 14654 5455 14688 5489
rect 15482 5455 15516 5489
rect 15554 5455 15588 5489
rect 16382 5455 16416 5489
rect 16454 5455 16488 5489
rect 17282 5455 17316 5489
rect 17354 5455 17388 5489
rect 18182 5455 18216 5489
rect 18254 5455 18288 5489
<< poly >>
rect 2024 8590 2424 8606
rect 2024 8556 2071 8590
rect 2105 8556 2139 8590
rect 2173 8556 2207 8590
rect 2241 8556 2275 8590
rect 2309 8556 2343 8590
rect 2377 8556 2424 8590
rect 2024 8509 2424 8556
rect 3024 8590 3424 8606
rect 3024 8556 3071 8590
rect 3105 8556 3139 8590
rect 3173 8556 3207 8590
rect 3241 8556 3275 8590
rect 3309 8556 3343 8590
rect 3377 8556 3424 8590
rect 3024 8509 3424 8556
rect 2024 8062 2424 8109
rect 2024 8028 2071 8062
rect 2105 8028 2139 8062
rect 2173 8028 2207 8062
rect 2241 8028 2275 8062
rect 2309 8028 2343 8062
rect 2377 8028 2424 8062
rect 2024 8012 2424 8028
rect 3024 8062 3424 8109
rect 3024 8028 3071 8062
rect 3105 8028 3139 8062
rect 3173 8028 3207 8062
rect 3241 8028 3275 8062
rect 3309 8028 3343 8062
rect 3377 8028 3424 8062
rect 3024 8012 3424 8028
rect 2024 7850 2424 7866
rect 2024 7816 2071 7850
rect 2105 7816 2139 7850
rect 2173 7816 2207 7850
rect 2241 7816 2275 7850
rect 2309 7816 2343 7850
rect 2377 7816 2424 7850
rect 2024 7769 2424 7816
rect 3024 7850 3424 7866
rect 3024 7816 3071 7850
rect 3105 7816 3139 7850
rect 3173 7816 3207 7850
rect 3241 7816 3275 7850
rect 3309 7816 3343 7850
rect 3377 7816 3424 7850
rect 3024 7769 3424 7816
rect 2024 7322 2424 7369
rect 2024 7288 2071 7322
rect 2105 7288 2139 7322
rect 2173 7288 2207 7322
rect 2241 7288 2275 7322
rect 2309 7288 2343 7322
rect 2377 7288 2424 7322
rect 2024 7272 2424 7288
rect 3024 7322 3424 7369
rect 3024 7288 3071 7322
rect 3105 7288 3139 7322
rect 3173 7288 3207 7322
rect 3241 7288 3275 7322
rect 3309 7288 3343 7322
rect 3377 7288 3424 7322
rect 3024 7272 3424 7288
rect 11742 6930 12142 6946
rect 11742 6896 11789 6930
rect 11823 6896 11857 6930
rect 11891 6896 11925 6930
rect 11959 6896 11993 6930
rect 12027 6896 12061 6930
rect 12095 6896 12142 6930
rect 11742 6849 12142 6896
rect 12642 6930 13042 6946
rect 12642 6896 12689 6930
rect 12723 6896 12757 6930
rect 12791 6896 12825 6930
rect 12859 6896 12893 6930
rect 12927 6896 12961 6930
rect 12995 6896 13042 6930
rect 12642 6849 13042 6896
rect 13542 6930 13942 6946
rect 13542 6896 13589 6930
rect 13623 6896 13657 6930
rect 13691 6896 13725 6930
rect 13759 6896 13793 6930
rect 13827 6896 13861 6930
rect 13895 6896 13942 6930
rect 13542 6849 13942 6896
rect 14442 6930 14842 6946
rect 14442 6896 14489 6930
rect 14523 6896 14557 6930
rect 14591 6896 14625 6930
rect 14659 6896 14693 6930
rect 14727 6896 14761 6930
rect 14795 6896 14842 6930
rect 14442 6849 14842 6896
rect 15342 6930 15742 6946
rect 15342 6896 15389 6930
rect 15423 6896 15457 6930
rect 15491 6896 15525 6930
rect 15559 6896 15593 6930
rect 15627 6896 15661 6930
rect 15695 6896 15742 6930
rect 15342 6849 15742 6896
rect 16242 6930 16642 6946
rect 16242 6896 16289 6930
rect 16323 6896 16357 6930
rect 16391 6896 16425 6930
rect 16459 6896 16493 6930
rect 16527 6896 16561 6930
rect 16595 6896 16642 6930
rect 16242 6849 16642 6896
rect 17142 6930 17542 6946
rect 17142 6896 17189 6930
rect 17223 6896 17257 6930
rect 17291 6896 17325 6930
rect 17359 6896 17393 6930
rect 17427 6896 17461 6930
rect 17495 6896 17542 6930
rect 17142 6849 17542 6896
rect 18042 6930 18442 6946
rect 18042 6896 18089 6930
rect 18123 6896 18157 6930
rect 18191 6896 18225 6930
rect 18259 6896 18293 6930
rect 18327 6896 18361 6930
rect 18395 6896 18442 6930
rect 18042 6849 18442 6896
rect 11742 6402 12142 6449
rect 11742 6368 11789 6402
rect 11823 6368 11857 6402
rect 11891 6368 11925 6402
rect 11959 6368 11993 6402
rect 12027 6368 12061 6402
rect 12095 6368 12142 6402
rect 11742 6352 12142 6368
rect 12642 6402 13042 6449
rect 12642 6368 12689 6402
rect 12723 6368 12757 6402
rect 12791 6368 12825 6402
rect 12859 6368 12893 6402
rect 12927 6368 12961 6402
rect 12995 6368 13042 6402
rect 12642 6352 13042 6368
rect 13542 6402 13942 6449
rect 13542 6368 13589 6402
rect 13623 6368 13657 6402
rect 13691 6368 13725 6402
rect 13759 6368 13793 6402
rect 13827 6368 13861 6402
rect 13895 6368 13942 6402
rect 13542 6352 13942 6368
rect 14442 6402 14842 6449
rect 14442 6368 14489 6402
rect 14523 6368 14557 6402
rect 14591 6368 14625 6402
rect 14659 6368 14693 6402
rect 14727 6368 14761 6402
rect 14795 6368 14842 6402
rect 14442 6352 14842 6368
rect 15342 6402 15742 6449
rect 15342 6368 15389 6402
rect 15423 6368 15457 6402
rect 15491 6368 15525 6402
rect 15559 6368 15593 6402
rect 15627 6368 15661 6402
rect 15695 6368 15742 6402
rect 15342 6352 15742 6368
rect 16242 6402 16642 6449
rect 16242 6368 16289 6402
rect 16323 6368 16357 6402
rect 16391 6368 16425 6402
rect 16459 6368 16493 6402
rect 16527 6368 16561 6402
rect 16595 6368 16642 6402
rect 16242 6352 16642 6368
rect 17142 6402 17542 6449
rect 17142 6368 17189 6402
rect 17223 6368 17257 6402
rect 17291 6368 17325 6402
rect 17359 6368 17393 6402
rect 17427 6368 17461 6402
rect 17495 6368 17542 6402
rect 17142 6352 17542 6368
rect 18042 6402 18442 6449
rect 18042 6368 18089 6402
rect 18123 6368 18157 6402
rect 18191 6368 18225 6402
rect 18259 6368 18293 6402
rect 18327 6368 18361 6402
rect 18395 6368 18442 6402
rect 18042 6352 18442 6368
rect 11742 6190 12142 6206
rect 11742 6156 11789 6190
rect 11823 6156 11857 6190
rect 11891 6156 11925 6190
rect 11959 6156 11993 6190
rect 12027 6156 12061 6190
rect 12095 6156 12142 6190
rect 11742 6109 12142 6156
rect 12642 6190 13042 6206
rect 12642 6156 12689 6190
rect 12723 6156 12757 6190
rect 12791 6156 12825 6190
rect 12859 6156 12893 6190
rect 12927 6156 12961 6190
rect 12995 6156 13042 6190
rect 12642 6109 13042 6156
rect 13542 6190 13942 6206
rect 13542 6156 13589 6190
rect 13623 6156 13657 6190
rect 13691 6156 13725 6190
rect 13759 6156 13793 6190
rect 13827 6156 13861 6190
rect 13895 6156 13942 6190
rect 13542 6109 13942 6156
rect 14442 6190 14842 6206
rect 14442 6156 14489 6190
rect 14523 6156 14557 6190
rect 14591 6156 14625 6190
rect 14659 6156 14693 6190
rect 14727 6156 14761 6190
rect 14795 6156 14842 6190
rect 14442 6109 14842 6156
rect 15342 6190 15742 6206
rect 15342 6156 15389 6190
rect 15423 6156 15457 6190
rect 15491 6156 15525 6190
rect 15559 6156 15593 6190
rect 15627 6156 15661 6190
rect 15695 6156 15742 6190
rect 15342 6109 15742 6156
rect 16242 6190 16642 6206
rect 16242 6156 16289 6190
rect 16323 6156 16357 6190
rect 16391 6156 16425 6190
rect 16459 6156 16493 6190
rect 16527 6156 16561 6190
rect 16595 6156 16642 6190
rect 16242 6109 16642 6156
rect 17142 6190 17542 6206
rect 17142 6156 17189 6190
rect 17223 6156 17257 6190
rect 17291 6156 17325 6190
rect 17359 6156 17393 6190
rect 17427 6156 17461 6190
rect 17495 6156 17542 6190
rect 17142 6109 17542 6156
rect 18042 6190 18442 6206
rect 18042 6156 18089 6190
rect 18123 6156 18157 6190
rect 18191 6156 18225 6190
rect 18259 6156 18293 6190
rect 18327 6156 18361 6190
rect 18395 6156 18442 6190
rect 18042 6109 18442 6156
rect -4208 5702 -4008 5718
rect -4208 5668 -4159 5702
rect -4125 5668 -4091 5702
rect -4057 5668 -4008 5702
rect -4208 5630 -4008 5668
rect -3508 5702 -3308 5718
rect -3508 5668 -3459 5702
rect -3425 5668 -3391 5702
rect -3357 5668 -3308 5702
rect -3508 5630 -3308 5668
rect -2808 5702 -2608 5718
rect -2808 5668 -2759 5702
rect -2725 5668 -2691 5702
rect -2657 5668 -2608 5702
rect -2808 5630 -2608 5668
rect -2108 5702 -1908 5718
rect -2108 5668 -2059 5702
rect -2025 5668 -1991 5702
rect -1957 5668 -1908 5702
rect -2108 5630 -1908 5668
rect -1408 5702 -1208 5718
rect -1408 5668 -1359 5702
rect -1325 5668 -1291 5702
rect -1257 5668 -1208 5702
rect -1408 5630 -1208 5668
rect -708 5702 -508 5718
rect -708 5668 -659 5702
rect -625 5668 -591 5702
rect -557 5668 -508 5702
rect -708 5630 -508 5668
rect -8 5702 192 5718
rect -8 5668 41 5702
rect 75 5668 109 5702
rect 143 5668 192 5702
rect -8 5630 192 5668
rect 692 5702 892 5718
rect 692 5668 741 5702
rect 775 5668 809 5702
rect 843 5668 892 5702
rect 692 5630 892 5668
rect 1392 5702 1592 5718
rect 1392 5668 1441 5702
rect 1475 5668 1509 5702
rect 1543 5668 1592 5702
rect 1392 5630 1592 5668
rect 2092 5702 2292 5718
rect 2092 5668 2141 5702
rect 2175 5668 2209 5702
rect 2243 5668 2292 5702
rect 2092 5630 2292 5668
rect 3792 5702 3992 5718
rect 3792 5668 3841 5702
rect 3875 5668 3909 5702
rect 3943 5668 3992 5702
rect 3792 5630 3992 5668
rect 4492 5702 4692 5718
rect 4492 5668 4541 5702
rect 4575 5668 4609 5702
rect 4643 5668 4692 5702
rect 4492 5630 4692 5668
rect 5192 5702 5392 5718
rect 5192 5668 5241 5702
rect 5275 5668 5309 5702
rect 5343 5668 5392 5702
rect 5192 5630 5392 5668
rect 5892 5702 6092 5718
rect 5892 5668 5941 5702
rect 5975 5668 6009 5702
rect 6043 5668 6092 5702
rect 5892 5630 6092 5668
rect 6592 5702 6792 5718
rect 6592 5668 6641 5702
rect 6675 5668 6709 5702
rect 6743 5668 6792 5702
rect 6592 5630 6792 5668
rect 7292 5702 7492 5718
rect 7292 5668 7341 5702
rect 7375 5668 7409 5702
rect 7443 5668 7492 5702
rect 7292 5630 7492 5668
rect 7992 5702 8192 5718
rect 7992 5668 8041 5702
rect 8075 5668 8109 5702
rect 8143 5668 8192 5702
rect 7992 5630 8192 5668
rect 8692 5702 8892 5718
rect 8692 5668 8741 5702
rect 8775 5668 8809 5702
rect 8843 5668 8892 5702
rect 8692 5630 8892 5668
rect 9392 5702 9592 5718
rect 9392 5668 9441 5702
rect 9475 5668 9509 5702
rect 9543 5668 9592 5702
rect 9392 5630 9592 5668
rect 10092 5702 10292 5718
rect 10092 5668 10141 5702
rect 10175 5668 10209 5702
rect 10243 5668 10292 5702
rect 10092 5630 10292 5668
rect 11742 5662 12142 5709
rect 11742 5628 11789 5662
rect 11823 5628 11857 5662
rect 11891 5628 11925 5662
rect 11959 5628 11993 5662
rect 12027 5628 12061 5662
rect 12095 5628 12142 5662
rect 11742 5612 12142 5628
rect 12642 5662 13042 5709
rect 12642 5628 12689 5662
rect 12723 5628 12757 5662
rect 12791 5628 12825 5662
rect 12859 5628 12893 5662
rect 12927 5628 12961 5662
rect 12995 5628 13042 5662
rect 12642 5612 13042 5628
rect 13542 5662 13942 5709
rect 13542 5628 13589 5662
rect 13623 5628 13657 5662
rect 13691 5628 13725 5662
rect 13759 5628 13793 5662
rect 13827 5628 13861 5662
rect 13895 5628 13942 5662
rect 13542 5612 13942 5628
rect 14442 5662 14842 5709
rect 14442 5628 14489 5662
rect 14523 5628 14557 5662
rect 14591 5628 14625 5662
rect 14659 5628 14693 5662
rect 14727 5628 14761 5662
rect 14795 5628 14842 5662
rect 14442 5612 14842 5628
rect 15342 5662 15742 5709
rect 15342 5628 15389 5662
rect 15423 5628 15457 5662
rect 15491 5628 15525 5662
rect 15559 5628 15593 5662
rect 15627 5628 15661 5662
rect 15695 5628 15742 5662
rect 15342 5612 15742 5628
rect 16242 5662 16642 5709
rect 16242 5628 16289 5662
rect 16323 5628 16357 5662
rect 16391 5628 16425 5662
rect 16459 5628 16493 5662
rect 16527 5628 16561 5662
rect 16595 5628 16642 5662
rect 16242 5612 16642 5628
rect 17142 5662 17542 5709
rect 17142 5628 17189 5662
rect 17223 5628 17257 5662
rect 17291 5628 17325 5662
rect 17359 5628 17393 5662
rect 17427 5628 17461 5662
rect 17495 5628 17542 5662
rect 17142 5612 17542 5628
rect 18042 5662 18442 5709
rect 18042 5628 18089 5662
rect 18123 5628 18157 5662
rect 18191 5628 18225 5662
rect 18259 5628 18293 5662
rect 18327 5628 18361 5662
rect 18395 5628 18442 5662
rect 18042 5612 18442 5628
rect -4208 3592 -4008 3630
rect -4208 3558 -4159 3592
rect -4125 3558 -4091 3592
rect -4057 3558 -4008 3592
rect -4208 3542 -4008 3558
rect -3508 3592 -3308 3630
rect -3508 3558 -3459 3592
rect -3425 3558 -3391 3592
rect -3357 3558 -3308 3592
rect -3508 3542 -3308 3558
rect -2808 3592 -2608 3630
rect -2808 3558 -2759 3592
rect -2725 3558 -2691 3592
rect -2657 3558 -2608 3592
rect -2808 3542 -2608 3558
rect -2108 3592 -1908 3630
rect -2108 3558 -2059 3592
rect -2025 3558 -1991 3592
rect -1957 3558 -1908 3592
rect -2108 3542 -1908 3558
rect -1408 3592 -1208 3630
rect -1408 3558 -1359 3592
rect -1325 3558 -1291 3592
rect -1257 3558 -1208 3592
rect -1408 3542 -1208 3558
rect -708 3592 -508 3630
rect -708 3558 -659 3592
rect -625 3558 -591 3592
rect -557 3558 -508 3592
rect -708 3542 -508 3558
rect -8 3592 192 3630
rect -8 3558 41 3592
rect 75 3558 109 3592
rect 143 3558 192 3592
rect -8 3542 192 3558
rect 692 3592 892 3630
rect 692 3558 741 3592
rect 775 3558 809 3592
rect 843 3558 892 3592
rect 692 3542 892 3558
rect 1392 3592 1592 3630
rect 1392 3558 1441 3592
rect 1475 3558 1509 3592
rect 1543 3558 1592 3592
rect 1392 3542 1592 3558
rect 2092 3592 2292 3630
rect 2092 3558 2141 3592
rect 2175 3558 2209 3592
rect 2243 3558 2292 3592
rect 2092 3542 2292 3558
rect 3792 3592 3992 3630
rect 3792 3558 3841 3592
rect 3875 3558 3909 3592
rect 3943 3558 3992 3592
rect 3792 3542 3992 3558
rect 4492 3592 4692 3630
rect 4492 3558 4541 3592
rect 4575 3558 4609 3592
rect 4643 3558 4692 3592
rect 4492 3542 4692 3558
rect 5192 3592 5392 3630
rect 5192 3558 5241 3592
rect 5275 3558 5309 3592
rect 5343 3558 5392 3592
rect 5192 3542 5392 3558
rect 5892 3592 6092 3630
rect 5892 3558 5941 3592
rect 5975 3558 6009 3592
rect 6043 3558 6092 3592
rect 5892 3542 6092 3558
rect 6592 3592 6792 3630
rect 6592 3558 6641 3592
rect 6675 3558 6709 3592
rect 6743 3558 6792 3592
rect 6592 3542 6792 3558
rect 7292 3592 7492 3630
rect 7292 3558 7341 3592
rect 7375 3558 7409 3592
rect 7443 3558 7492 3592
rect 7292 3542 7492 3558
rect 7992 3592 8192 3630
rect 7992 3558 8041 3592
rect 8075 3558 8109 3592
rect 8143 3558 8192 3592
rect 7992 3542 8192 3558
rect 8692 3592 8892 3630
rect 8692 3558 8741 3592
rect 8775 3558 8809 3592
rect 8843 3558 8892 3592
rect 8692 3542 8892 3558
rect 9392 3592 9592 3630
rect 9392 3558 9441 3592
rect 9475 3558 9509 3592
rect 9543 3558 9592 3592
rect 9392 3542 9592 3558
rect 10092 3592 10292 3630
rect 10092 3558 10141 3592
rect 10175 3558 10209 3592
rect 10243 3558 10292 3592
rect 10092 3542 10292 3558
rect 1134 1988 1534 2004
rect 1134 1954 1181 1988
rect 1215 1954 1249 1988
rect 1283 1954 1317 1988
rect 1351 1954 1385 1988
rect 1419 1954 1453 1988
rect 1487 1954 1534 1988
rect 1134 1916 1534 1954
rect 2134 1988 2534 2004
rect 2134 1954 2181 1988
rect 2215 1954 2249 1988
rect 2283 1954 2317 1988
rect 2351 1954 2385 1988
rect 2419 1954 2453 1988
rect 2487 1954 2534 1988
rect 2134 1916 2534 1954
rect 3134 1988 3534 2004
rect 3134 1954 3181 1988
rect 3215 1954 3249 1988
rect 3283 1954 3317 1988
rect 3351 1954 3385 1988
rect 3419 1954 3453 1988
rect 3487 1954 3534 1988
rect 3134 1916 3534 1954
rect 4134 1988 4534 2004
rect 4134 1954 4181 1988
rect 4215 1954 4249 1988
rect 4283 1954 4317 1988
rect 4351 1954 4385 1988
rect 4419 1954 4453 1988
rect 4487 1954 4534 1988
rect 4134 1916 4534 1954
rect 5134 1988 5534 2004
rect 5134 1954 5181 1988
rect 5215 1954 5249 1988
rect 5283 1954 5317 1988
rect 5351 1954 5385 1988
rect 5419 1954 5453 1988
rect 5487 1954 5534 1988
rect 5134 1916 5534 1954
rect 6134 1988 6534 2004
rect 6134 1954 6181 1988
rect 6215 1954 6249 1988
rect 6283 1954 6317 1988
rect 6351 1954 6385 1988
rect 6419 1954 6453 1988
rect 6487 1954 6534 1988
rect 6134 1916 6534 1954
rect 7134 1988 7534 2004
rect 7134 1954 7181 1988
rect 7215 1954 7249 1988
rect 7283 1954 7317 1988
rect 7351 1954 7385 1988
rect 7419 1954 7453 1988
rect 7487 1954 7534 1988
rect 7134 1916 7534 1954
rect 8134 1988 8534 2004
rect 8134 1954 8181 1988
rect 8215 1954 8249 1988
rect 8283 1954 8317 1988
rect 8351 1954 8385 1988
rect 8419 1954 8453 1988
rect 8487 1954 8534 1988
rect 8134 1916 8534 1954
rect 9134 1988 9534 2004
rect 9134 1954 9181 1988
rect 9215 1954 9249 1988
rect 9283 1954 9317 1988
rect 9351 1954 9385 1988
rect 9419 1954 9453 1988
rect 9487 1954 9534 1988
rect 9134 1916 9534 1954
rect 10134 1988 10534 2004
rect 10134 1954 10181 1988
rect 10215 1954 10249 1988
rect 10283 1954 10317 1988
rect 10351 1954 10385 1988
rect 10419 1954 10453 1988
rect 10487 1954 10534 1988
rect 10134 1916 10534 1954
rect 1134 1678 1534 1716
rect 1134 1644 1181 1678
rect 1215 1644 1249 1678
rect 1283 1644 1317 1678
rect 1351 1644 1385 1678
rect 1419 1644 1453 1678
rect 1487 1644 1534 1678
rect 1134 1628 1534 1644
rect 2134 1678 2534 1716
rect 2134 1644 2181 1678
rect 2215 1644 2249 1678
rect 2283 1644 2317 1678
rect 2351 1644 2385 1678
rect 2419 1644 2453 1678
rect 2487 1644 2534 1678
rect 2134 1628 2534 1644
rect 3134 1678 3534 1716
rect 3134 1644 3181 1678
rect 3215 1644 3249 1678
rect 3283 1644 3317 1678
rect 3351 1644 3385 1678
rect 3419 1644 3453 1678
rect 3487 1644 3534 1678
rect 3134 1628 3534 1644
rect 4134 1678 4534 1716
rect 4134 1644 4181 1678
rect 4215 1644 4249 1678
rect 4283 1644 4317 1678
rect 4351 1644 4385 1678
rect 4419 1644 4453 1678
rect 4487 1644 4534 1678
rect 4134 1628 4534 1644
rect 5134 1678 5534 1716
rect 5134 1644 5181 1678
rect 5215 1644 5249 1678
rect 5283 1644 5317 1678
rect 5351 1644 5385 1678
rect 5419 1644 5453 1678
rect 5487 1644 5534 1678
rect 5134 1628 5534 1644
rect 6134 1678 6534 1716
rect 6134 1644 6181 1678
rect 6215 1644 6249 1678
rect 6283 1644 6317 1678
rect 6351 1644 6385 1678
rect 6419 1644 6453 1678
rect 6487 1644 6534 1678
rect 6134 1628 6534 1644
rect 7134 1678 7534 1716
rect 7134 1644 7181 1678
rect 7215 1644 7249 1678
rect 7283 1644 7317 1678
rect 7351 1644 7385 1678
rect 7419 1644 7453 1678
rect 7487 1644 7534 1678
rect 7134 1628 7534 1644
rect 8134 1678 8534 1716
rect 8134 1644 8181 1678
rect 8215 1644 8249 1678
rect 8283 1644 8317 1678
rect 8351 1644 8385 1678
rect 8419 1644 8453 1678
rect 8487 1644 8534 1678
rect 8134 1628 8534 1644
rect 9134 1678 9534 1716
rect 9134 1644 9181 1678
rect 9215 1644 9249 1678
rect 9283 1644 9317 1678
rect 9351 1644 9385 1678
rect 9419 1644 9453 1678
rect 9487 1644 9534 1678
rect 9134 1628 9534 1644
rect 10134 1678 10534 1716
rect 10134 1644 10181 1678
rect 10215 1644 10249 1678
rect 10283 1644 10317 1678
rect 10351 1644 10385 1678
rect 10419 1644 10453 1678
rect 10487 1644 10534 1678
rect 10134 1628 10534 1644
rect 1134 1488 1534 1504
rect 1134 1454 1181 1488
rect 1215 1454 1249 1488
rect 1283 1454 1317 1488
rect 1351 1454 1385 1488
rect 1419 1454 1453 1488
rect 1487 1454 1534 1488
rect 1134 1416 1534 1454
rect 2134 1488 2534 1504
rect 2134 1454 2181 1488
rect 2215 1454 2249 1488
rect 2283 1454 2317 1488
rect 2351 1454 2385 1488
rect 2419 1454 2453 1488
rect 2487 1454 2534 1488
rect 2134 1416 2534 1454
rect 3134 1488 3534 1504
rect 3134 1454 3181 1488
rect 3215 1454 3249 1488
rect 3283 1454 3317 1488
rect 3351 1454 3385 1488
rect 3419 1454 3453 1488
rect 3487 1454 3534 1488
rect 3134 1416 3534 1454
rect 4134 1488 4534 1504
rect 4134 1454 4181 1488
rect 4215 1454 4249 1488
rect 4283 1454 4317 1488
rect 4351 1454 4385 1488
rect 4419 1454 4453 1488
rect 4487 1454 4534 1488
rect 4134 1416 4534 1454
rect 5134 1488 5534 1504
rect 5134 1454 5181 1488
rect 5215 1454 5249 1488
rect 5283 1454 5317 1488
rect 5351 1454 5385 1488
rect 5419 1454 5453 1488
rect 5487 1454 5534 1488
rect 5134 1416 5534 1454
rect 6134 1488 6534 1504
rect 6134 1454 6181 1488
rect 6215 1454 6249 1488
rect 6283 1454 6317 1488
rect 6351 1454 6385 1488
rect 6419 1454 6453 1488
rect 6487 1454 6534 1488
rect 6134 1416 6534 1454
rect 7134 1488 7534 1504
rect 7134 1454 7181 1488
rect 7215 1454 7249 1488
rect 7283 1454 7317 1488
rect 7351 1454 7385 1488
rect 7419 1454 7453 1488
rect 7487 1454 7534 1488
rect 7134 1416 7534 1454
rect 8134 1488 8534 1504
rect 8134 1454 8181 1488
rect 8215 1454 8249 1488
rect 8283 1454 8317 1488
rect 8351 1454 8385 1488
rect 8419 1454 8453 1488
rect 8487 1454 8534 1488
rect 8134 1416 8534 1454
rect 9134 1488 9534 1504
rect 9134 1454 9181 1488
rect 9215 1454 9249 1488
rect 9283 1454 9317 1488
rect 9351 1454 9385 1488
rect 9419 1454 9453 1488
rect 9487 1454 9534 1488
rect 9134 1416 9534 1454
rect 10134 1488 10534 1504
rect 10134 1454 10181 1488
rect 10215 1454 10249 1488
rect 10283 1454 10317 1488
rect 10351 1454 10385 1488
rect 10419 1454 10453 1488
rect 10487 1454 10534 1488
rect 10134 1416 10534 1454
rect 1134 1178 1534 1216
rect 1134 1144 1181 1178
rect 1215 1144 1249 1178
rect 1283 1144 1317 1178
rect 1351 1144 1385 1178
rect 1419 1144 1453 1178
rect 1487 1144 1534 1178
rect 1134 1128 1534 1144
rect 2134 1178 2534 1216
rect 2134 1144 2181 1178
rect 2215 1144 2249 1178
rect 2283 1144 2317 1178
rect 2351 1144 2385 1178
rect 2419 1144 2453 1178
rect 2487 1144 2534 1178
rect 2134 1128 2534 1144
rect 3134 1178 3534 1216
rect 3134 1144 3181 1178
rect 3215 1144 3249 1178
rect 3283 1144 3317 1178
rect 3351 1144 3385 1178
rect 3419 1144 3453 1178
rect 3487 1144 3534 1178
rect 3134 1128 3534 1144
rect 4134 1178 4534 1216
rect 4134 1144 4181 1178
rect 4215 1144 4249 1178
rect 4283 1144 4317 1178
rect 4351 1144 4385 1178
rect 4419 1144 4453 1178
rect 4487 1144 4534 1178
rect 4134 1128 4534 1144
rect 5134 1178 5534 1216
rect 5134 1144 5181 1178
rect 5215 1144 5249 1178
rect 5283 1144 5317 1178
rect 5351 1144 5385 1178
rect 5419 1144 5453 1178
rect 5487 1144 5534 1178
rect 5134 1128 5534 1144
rect 6134 1178 6534 1216
rect 6134 1144 6181 1178
rect 6215 1144 6249 1178
rect 6283 1144 6317 1178
rect 6351 1144 6385 1178
rect 6419 1144 6453 1178
rect 6487 1144 6534 1178
rect 6134 1128 6534 1144
rect 7134 1178 7534 1216
rect 7134 1144 7181 1178
rect 7215 1144 7249 1178
rect 7283 1144 7317 1178
rect 7351 1144 7385 1178
rect 7419 1144 7453 1178
rect 7487 1144 7534 1178
rect 7134 1128 7534 1144
rect 8134 1178 8534 1216
rect 8134 1144 8181 1178
rect 8215 1144 8249 1178
rect 8283 1144 8317 1178
rect 8351 1144 8385 1178
rect 8419 1144 8453 1178
rect 8487 1144 8534 1178
rect 8134 1128 8534 1144
rect 9134 1178 9534 1216
rect 9134 1144 9181 1178
rect 9215 1144 9249 1178
rect 9283 1144 9317 1178
rect 9351 1144 9385 1178
rect 9419 1144 9453 1178
rect 9487 1144 9534 1178
rect 9134 1128 9534 1144
rect 10134 1178 10534 1216
rect 10134 1144 10181 1178
rect 10215 1144 10249 1178
rect 10283 1144 10317 1178
rect 10351 1144 10385 1178
rect 10419 1144 10453 1178
rect 10487 1144 10534 1178
rect 10134 1128 10534 1144
<< polycont >>
rect 2071 8556 2105 8590
rect 2139 8556 2173 8590
rect 2207 8556 2241 8590
rect 2275 8556 2309 8590
rect 2343 8556 2377 8590
rect 3071 8556 3105 8590
rect 3139 8556 3173 8590
rect 3207 8556 3241 8590
rect 3275 8556 3309 8590
rect 3343 8556 3377 8590
rect 2071 8028 2105 8062
rect 2139 8028 2173 8062
rect 2207 8028 2241 8062
rect 2275 8028 2309 8062
rect 2343 8028 2377 8062
rect 3071 8028 3105 8062
rect 3139 8028 3173 8062
rect 3207 8028 3241 8062
rect 3275 8028 3309 8062
rect 3343 8028 3377 8062
rect 2071 7816 2105 7850
rect 2139 7816 2173 7850
rect 2207 7816 2241 7850
rect 2275 7816 2309 7850
rect 2343 7816 2377 7850
rect 3071 7816 3105 7850
rect 3139 7816 3173 7850
rect 3207 7816 3241 7850
rect 3275 7816 3309 7850
rect 3343 7816 3377 7850
rect 2071 7288 2105 7322
rect 2139 7288 2173 7322
rect 2207 7288 2241 7322
rect 2275 7288 2309 7322
rect 2343 7288 2377 7322
rect 3071 7288 3105 7322
rect 3139 7288 3173 7322
rect 3207 7288 3241 7322
rect 3275 7288 3309 7322
rect 3343 7288 3377 7322
rect 11789 6896 11823 6930
rect 11857 6896 11891 6930
rect 11925 6896 11959 6930
rect 11993 6896 12027 6930
rect 12061 6896 12095 6930
rect 12689 6896 12723 6930
rect 12757 6896 12791 6930
rect 12825 6896 12859 6930
rect 12893 6896 12927 6930
rect 12961 6896 12995 6930
rect 13589 6896 13623 6930
rect 13657 6896 13691 6930
rect 13725 6896 13759 6930
rect 13793 6896 13827 6930
rect 13861 6896 13895 6930
rect 14489 6896 14523 6930
rect 14557 6896 14591 6930
rect 14625 6896 14659 6930
rect 14693 6896 14727 6930
rect 14761 6896 14795 6930
rect 15389 6896 15423 6930
rect 15457 6896 15491 6930
rect 15525 6896 15559 6930
rect 15593 6896 15627 6930
rect 15661 6896 15695 6930
rect 16289 6896 16323 6930
rect 16357 6896 16391 6930
rect 16425 6896 16459 6930
rect 16493 6896 16527 6930
rect 16561 6896 16595 6930
rect 17189 6896 17223 6930
rect 17257 6896 17291 6930
rect 17325 6896 17359 6930
rect 17393 6896 17427 6930
rect 17461 6896 17495 6930
rect 18089 6896 18123 6930
rect 18157 6896 18191 6930
rect 18225 6896 18259 6930
rect 18293 6896 18327 6930
rect 18361 6896 18395 6930
rect 11789 6368 11823 6402
rect 11857 6368 11891 6402
rect 11925 6368 11959 6402
rect 11993 6368 12027 6402
rect 12061 6368 12095 6402
rect 12689 6368 12723 6402
rect 12757 6368 12791 6402
rect 12825 6368 12859 6402
rect 12893 6368 12927 6402
rect 12961 6368 12995 6402
rect 13589 6368 13623 6402
rect 13657 6368 13691 6402
rect 13725 6368 13759 6402
rect 13793 6368 13827 6402
rect 13861 6368 13895 6402
rect 14489 6368 14523 6402
rect 14557 6368 14591 6402
rect 14625 6368 14659 6402
rect 14693 6368 14727 6402
rect 14761 6368 14795 6402
rect 15389 6368 15423 6402
rect 15457 6368 15491 6402
rect 15525 6368 15559 6402
rect 15593 6368 15627 6402
rect 15661 6368 15695 6402
rect 16289 6368 16323 6402
rect 16357 6368 16391 6402
rect 16425 6368 16459 6402
rect 16493 6368 16527 6402
rect 16561 6368 16595 6402
rect 17189 6368 17223 6402
rect 17257 6368 17291 6402
rect 17325 6368 17359 6402
rect 17393 6368 17427 6402
rect 17461 6368 17495 6402
rect 18089 6368 18123 6402
rect 18157 6368 18191 6402
rect 18225 6368 18259 6402
rect 18293 6368 18327 6402
rect 18361 6368 18395 6402
rect 11789 6156 11823 6190
rect 11857 6156 11891 6190
rect 11925 6156 11959 6190
rect 11993 6156 12027 6190
rect 12061 6156 12095 6190
rect 12689 6156 12723 6190
rect 12757 6156 12791 6190
rect 12825 6156 12859 6190
rect 12893 6156 12927 6190
rect 12961 6156 12995 6190
rect 13589 6156 13623 6190
rect 13657 6156 13691 6190
rect 13725 6156 13759 6190
rect 13793 6156 13827 6190
rect 13861 6156 13895 6190
rect 14489 6156 14523 6190
rect 14557 6156 14591 6190
rect 14625 6156 14659 6190
rect 14693 6156 14727 6190
rect 14761 6156 14795 6190
rect 15389 6156 15423 6190
rect 15457 6156 15491 6190
rect 15525 6156 15559 6190
rect 15593 6156 15627 6190
rect 15661 6156 15695 6190
rect 16289 6156 16323 6190
rect 16357 6156 16391 6190
rect 16425 6156 16459 6190
rect 16493 6156 16527 6190
rect 16561 6156 16595 6190
rect 17189 6156 17223 6190
rect 17257 6156 17291 6190
rect 17325 6156 17359 6190
rect 17393 6156 17427 6190
rect 17461 6156 17495 6190
rect 18089 6156 18123 6190
rect 18157 6156 18191 6190
rect 18225 6156 18259 6190
rect 18293 6156 18327 6190
rect 18361 6156 18395 6190
rect -4159 5668 -4125 5702
rect -4091 5668 -4057 5702
rect -3459 5668 -3425 5702
rect -3391 5668 -3357 5702
rect -2759 5668 -2725 5702
rect -2691 5668 -2657 5702
rect -2059 5668 -2025 5702
rect -1991 5668 -1957 5702
rect -1359 5668 -1325 5702
rect -1291 5668 -1257 5702
rect -659 5668 -625 5702
rect -591 5668 -557 5702
rect 41 5668 75 5702
rect 109 5668 143 5702
rect 741 5668 775 5702
rect 809 5668 843 5702
rect 1441 5668 1475 5702
rect 1509 5668 1543 5702
rect 2141 5668 2175 5702
rect 2209 5668 2243 5702
rect 3841 5668 3875 5702
rect 3909 5668 3943 5702
rect 4541 5668 4575 5702
rect 4609 5668 4643 5702
rect 5241 5668 5275 5702
rect 5309 5668 5343 5702
rect 5941 5668 5975 5702
rect 6009 5668 6043 5702
rect 6641 5668 6675 5702
rect 6709 5668 6743 5702
rect 7341 5668 7375 5702
rect 7409 5668 7443 5702
rect 8041 5668 8075 5702
rect 8109 5668 8143 5702
rect 8741 5668 8775 5702
rect 8809 5668 8843 5702
rect 9441 5668 9475 5702
rect 9509 5668 9543 5702
rect 10141 5668 10175 5702
rect 10209 5668 10243 5702
rect 11789 5628 11823 5662
rect 11857 5628 11891 5662
rect 11925 5628 11959 5662
rect 11993 5628 12027 5662
rect 12061 5628 12095 5662
rect 12689 5628 12723 5662
rect 12757 5628 12791 5662
rect 12825 5628 12859 5662
rect 12893 5628 12927 5662
rect 12961 5628 12995 5662
rect 13589 5628 13623 5662
rect 13657 5628 13691 5662
rect 13725 5628 13759 5662
rect 13793 5628 13827 5662
rect 13861 5628 13895 5662
rect 14489 5628 14523 5662
rect 14557 5628 14591 5662
rect 14625 5628 14659 5662
rect 14693 5628 14727 5662
rect 14761 5628 14795 5662
rect 15389 5628 15423 5662
rect 15457 5628 15491 5662
rect 15525 5628 15559 5662
rect 15593 5628 15627 5662
rect 15661 5628 15695 5662
rect 16289 5628 16323 5662
rect 16357 5628 16391 5662
rect 16425 5628 16459 5662
rect 16493 5628 16527 5662
rect 16561 5628 16595 5662
rect 17189 5628 17223 5662
rect 17257 5628 17291 5662
rect 17325 5628 17359 5662
rect 17393 5628 17427 5662
rect 17461 5628 17495 5662
rect 18089 5628 18123 5662
rect 18157 5628 18191 5662
rect 18225 5628 18259 5662
rect 18293 5628 18327 5662
rect 18361 5628 18395 5662
rect -4159 3558 -4125 3592
rect -4091 3558 -4057 3592
rect -3459 3558 -3425 3592
rect -3391 3558 -3357 3592
rect -2759 3558 -2725 3592
rect -2691 3558 -2657 3592
rect -2059 3558 -2025 3592
rect -1991 3558 -1957 3592
rect -1359 3558 -1325 3592
rect -1291 3558 -1257 3592
rect -659 3558 -625 3592
rect -591 3558 -557 3592
rect 41 3558 75 3592
rect 109 3558 143 3592
rect 741 3558 775 3592
rect 809 3558 843 3592
rect 1441 3558 1475 3592
rect 1509 3558 1543 3592
rect 2141 3558 2175 3592
rect 2209 3558 2243 3592
rect 3841 3558 3875 3592
rect 3909 3558 3943 3592
rect 4541 3558 4575 3592
rect 4609 3558 4643 3592
rect 5241 3558 5275 3592
rect 5309 3558 5343 3592
rect 5941 3558 5975 3592
rect 6009 3558 6043 3592
rect 6641 3558 6675 3592
rect 6709 3558 6743 3592
rect 7341 3558 7375 3592
rect 7409 3558 7443 3592
rect 8041 3558 8075 3592
rect 8109 3558 8143 3592
rect 8741 3558 8775 3592
rect 8809 3558 8843 3592
rect 9441 3558 9475 3592
rect 9509 3558 9543 3592
rect 10141 3558 10175 3592
rect 10209 3558 10243 3592
rect 1181 1954 1215 1988
rect 1249 1954 1283 1988
rect 1317 1954 1351 1988
rect 1385 1954 1419 1988
rect 1453 1954 1487 1988
rect 2181 1954 2215 1988
rect 2249 1954 2283 1988
rect 2317 1954 2351 1988
rect 2385 1954 2419 1988
rect 2453 1954 2487 1988
rect 3181 1954 3215 1988
rect 3249 1954 3283 1988
rect 3317 1954 3351 1988
rect 3385 1954 3419 1988
rect 3453 1954 3487 1988
rect 4181 1954 4215 1988
rect 4249 1954 4283 1988
rect 4317 1954 4351 1988
rect 4385 1954 4419 1988
rect 4453 1954 4487 1988
rect 5181 1954 5215 1988
rect 5249 1954 5283 1988
rect 5317 1954 5351 1988
rect 5385 1954 5419 1988
rect 5453 1954 5487 1988
rect 6181 1954 6215 1988
rect 6249 1954 6283 1988
rect 6317 1954 6351 1988
rect 6385 1954 6419 1988
rect 6453 1954 6487 1988
rect 7181 1954 7215 1988
rect 7249 1954 7283 1988
rect 7317 1954 7351 1988
rect 7385 1954 7419 1988
rect 7453 1954 7487 1988
rect 8181 1954 8215 1988
rect 8249 1954 8283 1988
rect 8317 1954 8351 1988
rect 8385 1954 8419 1988
rect 8453 1954 8487 1988
rect 9181 1954 9215 1988
rect 9249 1954 9283 1988
rect 9317 1954 9351 1988
rect 9385 1954 9419 1988
rect 9453 1954 9487 1988
rect 10181 1954 10215 1988
rect 10249 1954 10283 1988
rect 10317 1954 10351 1988
rect 10385 1954 10419 1988
rect 10453 1954 10487 1988
rect 1181 1644 1215 1678
rect 1249 1644 1283 1678
rect 1317 1644 1351 1678
rect 1385 1644 1419 1678
rect 1453 1644 1487 1678
rect 2181 1644 2215 1678
rect 2249 1644 2283 1678
rect 2317 1644 2351 1678
rect 2385 1644 2419 1678
rect 2453 1644 2487 1678
rect 3181 1644 3215 1678
rect 3249 1644 3283 1678
rect 3317 1644 3351 1678
rect 3385 1644 3419 1678
rect 3453 1644 3487 1678
rect 4181 1644 4215 1678
rect 4249 1644 4283 1678
rect 4317 1644 4351 1678
rect 4385 1644 4419 1678
rect 4453 1644 4487 1678
rect 5181 1644 5215 1678
rect 5249 1644 5283 1678
rect 5317 1644 5351 1678
rect 5385 1644 5419 1678
rect 5453 1644 5487 1678
rect 6181 1644 6215 1678
rect 6249 1644 6283 1678
rect 6317 1644 6351 1678
rect 6385 1644 6419 1678
rect 6453 1644 6487 1678
rect 7181 1644 7215 1678
rect 7249 1644 7283 1678
rect 7317 1644 7351 1678
rect 7385 1644 7419 1678
rect 7453 1644 7487 1678
rect 8181 1644 8215 1678
rect 8249 1644 8283 1678
rect 8317 1644 8351 1678
rect 8385 1644 8419 1678
rect 8453 1644 8487 1678
rect 9181 1644 9215 1678
rect 9249 1644 9283 1678
rect 9317 1644 9351 1678
rect 9385 1644 9419 1678
rect 9453 1644 9487 1678
rect 10181 1644 10215 1678
rect 10249 1644 10283 1678
rect 10317 1644 10351 1678
rect 10385 1644 10419 1678
rect 10453 1644 10487 1678
rect 1181 1454 1215 1488
rect 1249 1454 1283 1488
rect 1317 1454 1351 1488
rect 1385 1454 1419 1488
rect 1453 1454 1487 1488
rect 2181 1454 2215 1488
rect 2249 1454 2283 1488
rect 2317 1454 2351 1488
rect 2385 1454 2419 1488
rect 2453 1454 2487 1488
rect 3181 1454 3215 1488
rect 3249 1454 3283 1488
rect 3317 1454 3351 1488
rect 3385 1454 3419 1488
rect 3453 1454 3487 1488
rect 4181 1454 4215 1488
rect 4249 1454 4283 1488
rect 4317 1454 4351 1488
rect 4385 1454 4419 1488
rect 4453 1454 4487 1488
rect 5181 1454 5215 1488
rect 5249 1454 5283 1488
rect 5317 1454 5351 1488
rect 5385 1454 5419 1488
rect 5453 1454 5487 1488
rect 6181 1454 6215 1488
rect 6249 1454 6283 1488
rect 6317 1454 6351 1488
rect 6385 1454 6419 1488
rect 6453 1454 6487 1488
rect 7181 1454 7215 1488
rect 7249 1454 7283 1488
rect 7317 1454 7351 1488
rect 7385 1454 7419 1488
rect 7453 1454 7487 1488
rect 8181 1454 8215 1488
rect 8249 1454 8283 1488
rect 8317 1454 8351 1488
rect 8385 1454 8419 1488
rect 8453 1454 8487 1488
rect 9181 1454 9215 1488
rect 9249 1454 9283 1488
rect 9317 1454 9351 1488
rect 9385 1454 9419 1488
rect 9453 1454 9487 1488
rect 10181 1454 10215 1488
rect 10249 1454 10283 1488
rect 10317 1454 10351 1488
rect 10385 1454 10419 1488
rect 10453 1454 10487 1488
rect 1181 1144 1215 1178
rect 1249 1144 1283 1178
rect 1317 1144 1351 1178
rect 1385 1144 1419 1178
rect 1453 1144 1487 1178
rect 2181 1144 2215 1178
rect 2249 1144 2283 1178
rect 2317 1144 2351 1178
rect 2385 1144 2419 1178
rect 2453 1144 2487 1178
rect 3181 1144 3215 1178
rect 3249 1144 3283 1178
rect 3317 1144 3351 1178
rect 3385 1144 3419 1178
rect 3453 1144 3487 1178
rect 4181 1144 4215 1178
rect 4249 1144 4283 1178
rect 4317 1144 4351 1178
rect 4385 1144 4419 1178
rect 4453 1144 4487 1178
rect 5181 1144 5215 1178
rect 5249 1144 5283 1178
rect 5317 1144 5351 1178
rect 5385 1144 5419 1178
rect 5453 1144 5487 1178
rect 6181 1144 6215 1178
rect 6249 1144 6283 1178
rect 6317 1144 6351 1178
rect 6385 1144 6419 1178
rect 6453 1144 6487 1178
rect 7181 1144 7215 1178
rect 7249 1144 7283 1178
rect 7317 1144 7351 1178
rect 7385 1144 7419 1178
rect 7453 1144 7487 1178
rect 8181 1144 8215 1178
rect 8249 1144 8283 1178
rect 8317 1144 8351 1178
rect 8385 1144 8419 1178
rect 8453 1144 8487 1178
rect 9181 1144 9215 1178
rect 9249 1144 9283 1178
rect 9317 1144 9351 1178
rect 9385 1144 9419 1178
rect 9453 1144 9487 1178
rect 10181 1144 10215 1178
rect 10249 1144 10283 1178
rect 10317 1144 10351 1178
rect 10385 1144 10419 1178
rect 10453 1144 10487 1178
<< xpolycontact >>
rect 21439 8488 21577 8920
rect 21439 6056 21577 6488
<< xpolyres >>
rect 21439 6488 21577 8488
<< locali >>
rect 2151 8754 2289 8770
rect 2151 8720 2167 8754
rect 2201 8720 2239 8754
rect 2273 8720 2289 8754
rect 2151 8704 2289 8720
rect 3151 8754 3289 8770
rect 3151 8720 3167 8754
rect 3201 8720 3239 8754
rect 3273 8720 3289 8754
rect 3151 8704 3289 8720
rect 2024 8556 2063 8590
rect 2105 8556 2135 8590
rect 2173 8556 2207 8590
rect 2241 8556 2275 8590
rect 2313 8556 2343 8590
rect 2385 8556 2424 8590
rect 3024 8556 3063 8590
rect 3105 8556 3135 8590
rect 3173 8556 3207 8590
rect 3241 8556 3275 8590
rect 3313 8556 3343 8590
rect 3385 8556 3424 8590
rect 1978 8496 2012 8513
rect 1978 8428 2012 8436
rect 1978 8360 2012 8364
rect 1978 8254 2012 8258
rect 1978 8182 2012 8190
rect 1978 8105 2012 8122
rect 2436 8496 2470 8513
rect 2436 8428 2470 8436
rect 2436 8360 2470 8364
rect 2436 8254 2470 8258
rect 2436 8182 2470 8190
rect 2436 8105 2470 8122
rect 2978 8496 3012 8513
rect 2978 8428 3012 8436
rect 2978 8360 3012 8364
rect 2978 8254 3012 8258
rect 2978 8182 3012 8190
rect 2978 8105 3012 8122
rect 3436 8496 3470 8513
rect 3436 8428 3470 8436
rect 3436 8360 3470 8364
rect 3436 8254 3470 8258
rect 3436 8182 3470 8190
rect 3436 8105 3470 8122
rect 2024 8028 2063 8062
rect 2105 8028 2135 8062
rect 2173 8028 2207 8062
rect 2241 8028 2275 8062
rect 2313 8028 2343 8062
rect 2385 8028 2424 8062
rect 3024 8028 3063 8062
rect 3105 8028 3135 8062
rect 3173 8028 3207 8062
rect 3241 8028 3275 8062
rect 3313 8028 3343 8062
rect 3385 8028 3424 8062
rect 2024 7816 2063 7850
rect 2105 7816 2135 7850
rect 2173 7816 2207 7850
rect 2241 7816 2275 7850
rect 2313 7816 2343 7850
rect 2385 7816 2424 7850
rect 3024 7816 3063 7850
rect 3105 7816 3135 7850
rect 3173 7816 3207 7850
rect 3241 7816 3275 7850
rect 3313 7816 3343 7850
rect 3385 7816 3424 7850
rect 1978 7756 2012 7773
rect 1978 7688 2012 7696
rect 1978 7620 2012 7624
rect 1978 7514 2012 7518
rect 1978 7442 2012 7450
rect 1978 7365 2012 7382
rect 2436 7756 2470 7773
rect 2436 7688 2470 7696
rect 2436 7620 2470 7624
rect 2436 7514 2470 7518
rect 2436 7442 2470 7450
rect 2436 7365 2470 7382
rect 2978 7756 3012 7773
rect 2978 7688 3012 7696
rect 2978 7620 3012 7624
rect 2978 7514 3012 7518
rect 2978 7442 3012 7450
rect 2978 7365 3012 7382
rect 3436 7756 3470 7773
rect 3436 7688 3470 7696
rect 3436 7620 3470 7624
rect 3436 7514 3470 7518
rect 21081 7603 21147 7619
rect 21081 7568 21097 7603
rect 21131 7568 21147 7603
rect 21081 7531 21147 7568
rect 21081 7496 21097 7531
rect 21131 7496 21147 7531
rect 21081 7480 21147 7496
rect 3436 7442 3470 7450
rect 3436 7365 3470 7382
rect 2024 7288 2063 7322
rect 2105 7288 2135 7322
rect 2173 7288 2207 7322
rect 2241 7288 2275 7322
rect 2313 7288 2343 7322
rect 2385 7288 2424 7322
rect 3024 7288 3063 7322
rect 3105 7288 3135 7322
rect 3173 7288 3207 7322
rect 3241 7288 3275 7322
rect 3313 7288 3343 7322
rect 3385 7288 3424 7322
rect 2148 7149 2286 7165
rect 2148 7115 2164 7149
rect 2198 7115 2236 7149
rect 2270 7115 2286 7149
rect 2148 7099 2286 7115
rect 3148 7149 3286 7165
rect 3148 7115 3164 7149
rect 3198 7115 3236 7149
rect 3270 7115 3286 7149
rect 3148 7099 3286 7115
rect 11869 7094 12007 7110
rect 11869 7060 11885 7094
rect 11919 7060 11957 7094
rect 11991 7060 12007 7094
rect 11869 7044 12007 7060
rect 12769 7094 12907 7110
rect 12769 7060 12785 7094
rect 12819 7060 12857 7094
rect 12891 7060 12907 7094
rect 12769 7044 12907 7060
rect 13669 7094 13807 7110
rect 13669 7060 13685 7094
rect 13719 7060 13757 7094
rect 13791 7060 13807 7094
rect 13669 7044 13807 7060
rect 14569 7094 14707 7110
rect 14569 7060 14585 7094
rect 14619 7060 14657 7094
rect 14691 7060 14707 7094
rect 14569 7044 14707 7060
rect 15469 7094 15607 7110
rect 15469 7060 15485 7094
rect 15519 7060 15557 7094
rect 15591 7060 15607 7094
rect 15469 7044 15607 7060
rect 16369 7094 16507 7110
rect 16369 7060 16385 7094
rect 16419 7060 16457 7094
rect 16491 7060 16507 7094
rect 16369 7044 16507 7060
rect 17269 7094 17407 7110
rect 17269 7060 17285 7094
rect 17319 7060 17357 7094
rect 17391 7060 17407 7094
rect 17269 7044 17407 7060
rect 18169 7094 18307 7110
rect 18169 7060 18185 7094
rect 18219 7060 18257 7094
rect 18291 7060 18307 7094
rect 18169 7044 18307 7060
rect 11742 6896 11781 6930
rect 11823 6896 11853 6930
rect 11891 6896 11925 6930
rect 11959 6896 11993 6930
rect 12031 6896 12061 6930
rect 12103 6896 12142 6930
rect 12642 6896 12681 6930
rect 12723 6896 12753 6930
rect 12791 6896 12825 6930
rect 12859 6896 12893 6930
rect 12931 6896 12961 6930
rect 13003 6896 13042 6930
rect 13542 6896 13581 6930
rect 13623 6896 13653 6930
rect 13691 6896 13725 6930
rect 13759 6896 13793 6930
rect 13831 6896 13861 6930
rect 13903 6896 13942 6930
rect 14442 6896 14481 6930
rect 14523 6896 14553 6930
rect 14591 6896 14625 6930
rect 14659 6896 14693 6930
rect 14731 6896 14761 6930
rect 14803 6896 14842 6930
rect 15342 6896 15381 6930
rect 15423 6896 15453 6930
rect 15491 6896 15525 6930
rect 15559 6896 15593 6930
rect 15631 6896 15661 6930
rect 15703 6896 15742 6930
rect 16242 6896 16281 6930
rect 16323 6896 16353 6930
rect 16391 6896 16425 6930
rect 16459 6896 16493 6930
rect 16531 6896 16561 6930
rect 16603 6896 16642 6930
rect 17142 6896 17181 6930
rect 17223 6896 17253 6930
rect 17291 6896 17325 6930
rect 17359 6896 17393 6930
rect 17431 6896 17461 6930
rect 17503 6896 17542 6930
rect 18042 6896 18081 6930
rect 18123 6896 18153 6930
rect 18191 6896 18225 6930
rect 18259 6896 18293 6930
rect 18331 6896 18361 6930
rect 18403 6896 18442 6930
rect 11696 6836 11730 6853
rect 11696 6768 11730 6776
rect 11696 6700 11730 6704
rect 11696 6594 11730 6598
rect 11696 6522 11730 6530
rect 11696 6445 11730 6462
rect 12154 6836 12188 6853
rect 12154 6768 12188 6776
rect 12154 6700 12188 6704
rect 12154 6594 12188 6598
rect 12154 6522 12188 6530
rect 12154 6445 12188 6462
rect 12596 6836 12630 6853
rect 12596 6768 12630 6776
rect 12596 6700 12630 6704
rect 12596 6594 12630 6598
rect 12596 6522 12630 6530
rect 12596 6445 12630 6462
rect 13054 6836 13088 6853
rect 13054 6768 13088 6776
rect 13054 6700 13088 6704
rect 13054 6594 13088 6598
rect 13054 6522 13088 6530
rect 13054 6445 13088 6462
rect 13496 6836 13530 6853
rect 13496 6768 13530 6776
rect 13496 6700 13530 6704
rect 13496 6594 13530 6598
rect 13496 6522 13530 6530
rect 13496 6445 13530 6462
rect 13954 6836 13988 6853
rect 13954 6768 13988 6776
rect 13954 6700 13988 6704
rect 13954 6594 13988 6598
rect 13954 6522 13988 6530
rect 13954 6445 13988 6462
rect 14396 6836 14430 6853
rect 14396 6768 14430 6776
rect 14396 6700 14430 6704
rect 14396 6594 14430 6598
rect 14396 6522 14430 6530
rect 14396 6445 14430 6462
rect 14854 6836 14888 6853
rect 14854 6768 14888 6776
rect 14854 6700 14888 6704
rect 14854 6594 14888 6598
rect 14854 6522 14888 6530
rect 14854 6445 14888 6462
rect 15296 6836 15330 6853
rect 15296 6768 15330 6776
rect 15296 6700 15330 6704
rect 15296 6594 15330 6598
rect 15296 6522 15330 6530
rect 15296 6445 15330 6462
rect 15754 6836 15788 6853
rect 15754 6768 15788 6776
rect 15754 6700 15788 6704
rect 15754 6594 15788 6598
rect 15754 6522 15788 6530
rect 15754 6445 15788 6462
rect 16196 6836 16230 6853
rect 16196 6768 16230 6776
rect 16196 6700 16230 6704
rect 16196 6594 16230 6598
rect 16196 6522 16230 6530
rect 16196 6445 16230 6462
rect 16654 6836 16688 6853
rect 16654 6768 16688 6776
rect 16654 6700 16688 6704
rect 16654 6594 16688 6598
rect 16654 6522 16688 6530
rect 16654 6445 16688 6462
rect 17096 6836 17130 6853
rect 17096 6768 17130 6776
rect 17096 6700 17130 6704
rect 17096 6594 17130 6598
rect 17096 6522 17130 6530
rect 17096 6445 17130 6462
rect 17554 6836 17588 6853
rect 17554 6768 17588 6776
rect 17554 6700 17588 6704
rect 17554 6594 17588 6598
rect 17554 6522 17588 6530
rect 17554 6445 17588 6462
rect 17996 6836 18030 6853
rect 17996 6768 18030 6776
rect 17996 6700 18030 6704
rect 17996 6594 18030 6598
rect 17996 6522 18030 6530
rect 17996 6445 18030 6462
rect 18454 6836 18488 6853
rect 18454 6768 18488 6776
rect 18454 6700 18488 6704
rect 18454 6594 18488 6598
rect 18454 6522 18488 6530
rect 18454 6445 18488 6462
rect 11742 6368 11781 6402
rect 11823 6368 11853 6402
rect 11891 6368 11925 6402
rect 11959 6368 11993 6402
rect 12031 6368 12061 6402
rect 12103 6368 12142 6402
rect 12642 6368 12681 6402
rect 12723 6368 12753 6402
rect 12791 6368 12825 6402
rect 12859 6368 12893 6402
rect 12931 6368 12961 6402
rect 13003 6368 13042 6402
rect 13542 6368 13581 6402
rect 13623 6368 13653 6402
rect 13691 6368 13725 6402
rect 13759 6368 13793 6402
rect 13831 6368 13861 6402
rect 13903 6368 13942 6402
rect 14442 6368 14481 6402
rect 14523 6368 14553 6402
rect 14591 6368 14625 6402
rect 14659 6368 14693 6402
rect 14731 6368 14761 6402
rect 14803 6368 14842 6402
rect 15342 6368 15381 6402
rect 15423 6368 15453 6402
rect 15491 6368 15525 6402
rect 15559 6368 15593 6402
rect 15631 6368 15661 6402
rect 15703 6368 15742 6402
rect 16242 6368 16281 6402
rect 16323 6368 16353 6402
rect 16391 6368 16425 6402
rect 16459 6368 16493 6402
rect 16531 6368 16561 6402
rect 16603 6368 16642 6402
rect 17142 6368 17181 6402
rect 17223 6368 17253 6402
rect 17291 6368 17325 6402
rect 17359 6368 17393 6402
rect 17431 6368 17461 6402
rect 17503 6368 17542 6402
rect 18042 6368 18081 6402
rect 18123 6368 18153 6402
rect 18191 6368 18225 6402
rect 18259 6368 18293 6402
rect 18331 6368 18361 6402
rect 18403 6368 18442 6402
rect 11742 6156 11781 6190
rect 11823 6156 11853 6190
rect 11891 6156 11925 6190
rect 11959 6156 11993 6190
rect 12031 6156 12061 6190
rect 12103 6156 12142 6190
rect 12642 6156 12681 6190
rect 12723 6156 12753 6190
rect 12791 6156 12825 6190
rect 12859 6156 12893 6190
rect 12931 6156 12961 6190
rect 13003 6156 13042 6190
rect 13542 6156 13581 6190
rect 13623 6156 13653 6190
rect 13691 6156 13725 6190
rect 13759 6156 13793 6190
rect 13831 6156 13861 6190
rect 13903 6156 13942 6190
rect 14442 6156 14481 6190
rect 14523 6156 14553 6190
rect 14591 6156 14625 6190
rect 14659 6156 14693 6190
rect 14731 6156 14761 6190
rect 14803 6156 14842 6190
rect 15342 6156 15381 6190
rect 15423 6156 15453 6190
rect 15491 6156 15525 6190
rect 15559 6156 15593 6190
rect 15631 6156 15661 6190
rect 15703 6156 15742 6190
rect 16242 6156 16281 6190
rect 16323 6156 16353 6190
rect 16391 6156 16425 6190
rect 16459 6156 16493 6190
rect 16531 6156 16561 6190
rect 16603 6156 16642 6190
rect 17142 6156 17181 6190
rect 17223 6156 17253 6190
rect 17291 6156 17325 6190
rect 17359 6156 17393 6190
rect 17431 6156 17461 6190
rect 17503 6156 17542 6190
rect 18042 6156 18081 6190
rect 18123 6156 18153 6190
rect 18191 6156 18225 6190
rect 18259 6156 18293 6190
rect 18331 6156 18361 6190
rect 18403 6156 18442 6190
rect 11696 6096 11730 6113
rect 11696 6028 11730 6036
rect 11696 5960 11730 5964
rect -4168 5925 -4030 5941
rect -4168 5891 -4152 5925
rect -4118 5891 -4080 5925
rect -4046 5891 -4030 5925
rect -4168 5875 -4030 5891
rect -3468 5925 -3330 5941
rect -3468 5891 -3452 5925
rect -3418 5891 -3380 5925
rect -3346 5891 -3330 5925
rect -3468 5875 -3330 5891
rect -2768 5925 -2630 5941
rect -2768 5891 -2752 5925
rect -2718 5891 -2680 5925
rect -2646 5891 -2630 5925
rect -2768 5875 -2630 5891
rect -2068 5925 -1930 5941
rect -2068 5891 -2052 5925
rect -2018 5891 -1980 5925
rect -1946 5891 -1930 5925
rect -2068 5875 -1930 5891
rect -1368 5925 -1230 5941
rect -1368 5891 -1352 5925
rect -1318 5891 -1280 5925
rect -1246 5891 -1230 5925
rect -1368 5875 -1230 5891
rect -668 5925 -530 5941
rect -668 5891 -652 5925
rect -618 5891 -580 5925
rect -546 5891 -530 5925
rect -668 5875 -530 5891
rect 32 5925 170 5941
rect 32 5891 48 5925
rect 82 5891 120 5925
rect 154 5891 170 5925
rect 32 5875 170 5891
rect 732 5925 870 5941
rect 732 5891 748 5925
rect 782 5891 820 5925
rect 854 5891 870 5925
rect 732 5875 870 5891
rect 1432 5925 1570 5941
rect 1432 5891 1448 5925
rect 1482 5891 1520 5925
rect 1554 5891 1570 5925
rect 1432 5875 1570 5891
rect 2132 5925 2270 5941
rect 2132 5891 2148 5925
rect 2182 5891 2220 5925
rect 2254 5891 2270 5925
rect 2132 5875 2270 5891
rect 3832 5925 3970 5941
rect 3832 5891 3848 5925
rect 3882 5891 3920 5925
rect 3954 5891 3970 5925
rect 3832 5875 3970 5891
rect 4532 5925 4670 5941
rect 4532 5891 4548 5925
rect 4582 5891 4620 5925
rect 4654 5891 4670 5925
rect 4532 5875 4670 5891
rect 5232 5925 5370 5941
rect 5232 5891 5248 5925
rect 5282 5891 5320 5925
rect 5354 5891 5370 5925
rect 5232 5875 5370 5891
rect 5932 5925 6070 5941
rect 5932 5891 5948 5925
rect 5982 5891 6020 5925
rect 6054 5891 6070 5925
rect 5932 5875 6070 5891
rect 6632 5925 6770 5941
rect 6632 5891 6648 5925
rect 6682 5891 6720 5925
rect 6754 5891 6770 5925
rect 6632 5875 6770 5891
rect 7332 5925 7470 5941
rect 7332 5891 7348 5925
rect 7382 5891 7420 5925
rect 7454 5891 7470 5925
rect 7332 5875 7470 5891
rect 8032 5925 8170 5941
rect 8032 5891 8048 5925
rect 8082 5891 8120 5925
rect 8154 5891 8170 5925
rect 8032 5875 8170 5891
rect 8732 5925 8870 5941
rect 8732 5891 8748 5925
rect 8782 5891 8820 5925
rect 8854 5891 8870 5925
rect 8732 5875 8870 5891
rect 9432 5925 9570 5941
rect 9432 5891 9448 5925
rect 9482 5891 9520 5925
rect 9554 5891 9570 5925
rect 9432 5875 9570 5891
rect 10132 5925 10270 5941
rect 10132 5891 10148 5925
rect 10182 5891 10220 5925
rect 10254 5891 10270 5925
rect 10132 5875 10270 5891
rect 11696 5854 11730 5858
rect 11696 5782 11730 5790
rect 11696 5705 11730 5722
rect 12154 6096 12188 6113
rect 12154 6028 12188 6036
rect 12154 5960 12188 5964
rect 12154 5854 12188 5858
rect 12154 5782 12188 5790
rect 12154 5705 12188 5722
rect 12596 6096 12630 6113
rect 12596 6028 12630 6036
rect 12596 5960 12630 5964
rect 12596 5854 12630 5858
rect 12596 5782 12630 5790
rect 12596 5705 12630 5722
rect 13054 6096 13088 6113
rect 13054 6028 13088 6036
rect 13054 5960 13088 5964
rect 13054 5854 13088 5858
rect 13054 5782 13088 5790
rect 13054 5705 13088 5722
rect 13496 6096 13530 6113
rect 13496 6028 13530 6036
rect 13496 5960 13530 5964
rect 13496 5854 13530 5858
rect 13496 5782 13530 5790
rect 13496 5705 13530 5722
rect 13954 6096 13988 6113
rect 13954 6028 13988 6036
rect 13954 5960 13988 5964
rect 13954 5854 13988 5858
rect 13954 5782 13988 5790
rect 13954 5705 13988 5722
rect 14396 6096 14430 6113
rect 14396 6028 14430 6036
rect 14396 5960 14430 5964
rect 14396 5854 14430 5858
rect 14396 5782 14430 5790
rect 14396 5705 14430 5722
rect 14854 6096 14888 6113
rect 14854 6028 14888 6036
rect 14854 5960 14888 5964
rect 14854 5854 14888 5858
rect 14854 5782 14888 5790
rect 14854 5705 14888 5722
rect 15296 6096 15330 6113
rect 15296 6028 15330 6036
rect 15296 5960 15330 5964
rect 15296 5854 15330 5858
rect 15296 5782 15330 5790
rect 15296 5705 15330 5722
rect 15754 6096 15788 6113
rect 15754 6028 15788 6036
rect 15754 5960 15788 5964
rect 15754 5854 15788 5858
rect 15754 5782 15788 5790
rect 15754 5705 15788 5722
rect 16196 6096 16230 6113
rect 16196 6028 16230 6036
rect 16196 5960 16230 5964
rect 16196 5854 16230 5858
rect 16196 5782 16230 5790
rect 16196 5705 16230 5722
rect 16654 6096 16688 6113
rect 16654 6028 16688 6036
rect 16654 5960 16688 5964
rect 16654 5854 16688 5858
rect 16654 5782 16688 5790
rect 16654 5705 16688 5722
rect 17096 6096 17130 6113
rect 17096 6028 17130 6036
rect 17096 5960 17130 5964
rect 17096 5854 17130 5858
rect 17096 5782 17130 5790
rect 17096 5705 17130 5722
rect 17554 6096 17588 6113
rect 17554 6028 17588 6036
rect 17554 5960 17588 5964
rect 17554 5854 17588 5858
rect 17554 5782 17588 5790
rect 17554 5705 17588 5722
rect 17996 6096 18030 6113
rect 17996 6028 18030 6036
rect 17996 5960 18030 5964
rect 17996 5854 18030 5858
rect 17996 5782 18030 5790
rect 17996 5705 18030 5722
rect 18454 6096 18488 6113
rect 18454 6028 18488 6036
rect 18454 5960 18488 5964
rect 18454 5854 18488 5858
rect 18454 5782 18488 5790
rect 18454 5705 18488 5722
rect -4208 5668 -4161 5702
rect -4125 5668 -4091 5702
rect -4055 5668 -4008 5702
rect -3508 5668 -3461 5702
rect -3425 5668 -3391 5702
rect -3355 5668 -3308 5702
rect -2808 5668 -2761 5702
rect -2725 5668 -2691 5702
rect -2655 5668 -2608 5702
rect -2108 5668 -2061 5702
rect -2025 5668 -1991 5702
rect -1955 5668 -1908 5702
rect -1408 5668 -1361 5702
rect -1325 5668 -1291 5702
rect -1255 5668 -1208 5702
rect -708 5668 -661 5702
rect -625 5668 -591 5702
rect -555 5668 -508 5702
rect -8 5668 39 5702
rect 75 5668 109 5702
rect 145 5668 192 5702
rect 692 5668 739 5702
rect 775 5668 809 5702
rect 845 5668 892 5702
rect 1392 5668 1439 5702
rect 1475 5668 1509 5702
rect 1545 5668 1592 5702
rect 2092 5668 2139 5702
rect 2175 5668 2209 5702
rect 2245 5668 2292 5702
rect 3792 5668 3839 5702
rect 3875 5668 3909 5702
rect 3945 5668 3992 5702
rect 4492 5668 4539 5702
rect 4575 5668 4609 5702
rect 4645 5668 4692 5702
rect 5192 5668 5239 5702
rect 5275 5668 5309 5702
rect 5345 5668 5392 5702
rect 5892 5668 5939 5702
rect 5975 5668 6009 5702
rect 6045 5668 6092 5702
rect 6592 5668 6639 5702
rect 6675 5668 6709 5702
rect 6745 5668 6792 5702
rect 7292 5668 7339 5702
rect 7375 5668 7409 5702
rect 7445 5668 7492 5702
rect 7992 5668 8039 5702
rect 8075 5668 8109 5702
rect 8145 5668 8192 5702
rect 8692 5668 8739 5702
rect 8775 5668 8809 5702
rect 8845 5668 8892 5702
rect 9392 5668 9439 5702
rect 9475 5668 9509 5702
rect 9545 5668 9592 5702
rect 10092 5668 10139 5702
rect 10175 5668 10209 5702
rect 10245 5668 10292 5702
rect -4254 5599 -4220 5634
rect -4254 5531 -4220 5549
rect -4254 5463 -4220 5477
rect -4254 5395 -4220 5405
rect -4254 5327 -4220 5333
rect -4254 5259 -4220 5261
rect -4254 5223 -4220 5225
rect -4254 5151 -4220 5157
rect -4254 5079 -4220 5089
rect -4254 5007 -4220 5021
rect -4254 4935 -4220 4953
rect -4254 4863 -4220 4885
rect -4254 4791 -4220 4817
rect -4254 4719 -4220 4749
rect -4254 4647 -4220 4681
rect -4254 4579 -4220 4613
rect -4254 4511 -4220 4541
rect -4254 4443 -4220 4469
rect -4254 4375 -4220 4397
rect -4254 4307 -4220 4325
rect -4254 4239 -4220 4253
rect -4254 4171 -4220 4181
rect -4254 4103 -4220 4109
rect -4254 4035 -4220 4037
rect -4254 3999 -4220 4001
rect -4254 3927 -4220 3933
rect -4254 3855 -4220 3865
rect -4254 3783 -4220 3797
rect -4254 3711 -4220 3729
rect -4254 3626 -4220 3661
rect -3996 5599 -3962 5634
rect -3996 5531 -3962 5549
rect -3996 5463 -3962 5477
rect -3996 5395 -3962 5405
rect -3996 5327 -3962 5333
rect -3996 5259 -3962 5261
rect -3996 5223 -3962 5225
rect -3996 5151 -3962 5157
rect -3996 5079 -3962 5089
rect -3996 5007 -3962 5021
rect -3996 4935 -3962 4953
rect -3996 4863 -3962 4885
rect -3996 4791 -3962 4817
rect -3996 4719 -3962 4749
rect -3996 4647 -3962 4681
rect -3996 4579 -3962 4613
rect -3996 4511 -3962 4541
rect -3996 4443 -3962 4469
rect -3996 4375 -3962 4397
rect -3996 4307 -3962 4325
rect -3996 4239 -3962 4253
rect -3996 4171 -3962 4181
rect -3996 4103 -3962 4109
rect -3996 4035 -3962 4037
rect -3996 3999 -3962 4001
rect -3996 3927 -3962 3933
rect -3996 3855 -3962 3865
rect -3996 3783 -3962 3797
rect -3996 3711 -3962 3729
rect -3996 3626 -3962 3661
rect -3554 5599 -3520 5634
rect -3554 5531 -3520 5549
rect -3554 5463 -3520 5477
rect -3554 5395 -3520 5405
rect -3554 5327 -3520 5333
rect -3554 5259 -3520 5261
rect -3554 5223 -3520 5225
rect -3554 5151 -3520 5157
rect -3554 5079 -3520 5089
rect -3554 5007 -3520 5021
rect -3554 4935 -3520 4953
rect -3554 4863 -3520 4885
rect -3554 4791 -3520 4817
rect -3554 4719 -3520 4749
rect -3554 4647 -3520 4681
rect -3554 4579 -3520 4613
rect -3554 4511 -3520 4541
rect -3554 4443 -3520 4469
rect -3554 4375 -3520 4397
rect -3554 4307 -3520 4325
rect -3554 4239 -3520 4253
rect -3554 4171 -3520 4181
rect -3554 4103 -3520 4109
rect -3554 4035 -3520 4037
rect -3554 3999 -3520 4001
rect -3554 3927 -3520 3933
rect -3554 3855 -3520 3865
rect -3554 3783 -3520 3797
rect -3554 3711 -3520 3729
rect -3554 3626 -3520 3661
rect -3296 5599 -3262 5634
rect -3296 5531 -3262 5549
rect -3296 5463 -3262 5477
rect -3296 5395 -3262 5405
rect -3296 5327 -3262 5333
rect -3296 5259 -3262 5261
rect -3296 5223 -3262 5225
rect -3296 5151 -3262 5157
rect -3296 5079 -3262 5089
rect -3296 5007 -3262 5021
rect -3296 4935 -3262 4953
rect -3296 4863 -3262 4885
rect -3296 4791 -3262 4817
rect -3296 4719 -3262 4749
rect -3296 4647 -3262 4681
rect -3296 4579 -3262 4613
rect -3296 4511 -3262 4541
rect -3296 4443 -3262 4469
rect -3296 4375 -3262 4397
rect -3296 4307 -3262 4325
rect -3296 4239 -3262 4253
rect -3296 4171 -3262 4181
rect -3296 4103 -3262 4109
rect -3296 4035 -3262 4037
rect -3296 3999 -3262 4001
rect -3296 3927 -3262 3933
rect -3296 3855 -3262 3865
rect -3296 3783 -3262 3797
rect -3296 3711 -3262 3729
rect -3296 3626 -3262 3661
rect -2854 5599 -2820 5634
rect -2854 5531 -2820 5549
rect -2854 5463 -2820 5477
rect -2854 5395 -2820 5405
rect -2854 5327 -2820 5333
rect -2854 5259 -2820 5261
rect -2854 5223 -2820 5225
rect -2854 5151 -2820 5157
rect -2854 5079 -2820 5089
rect -2854 5007 -2820 5021
rect -2854 4935 -2820 4953
rect -2854 4863 -2820 4885
rect -2854 4791 -2820 4817
rect -2854 4719 -2820 4749
rect -2854 4647 -2820 4681
rect -2854 4579 -2820 4613
rect -2854 4511 -2820 4541
rect -2854 4443 -2820 4469
rect -2854 4375 -2820 4397
rect -2854 4307 -2820 4325
rect -2854 4239 -2820 4253
rect -2854 4171 -2820 4181
rect -2854 4103 -2820 4109
rect -2854 4035 -2820 4037
rect -2854 3999 -2820 4001
rect -2854 3927 -2820 3933
rect -2854 3855 -2820 3865
rect -2854 3783 -2820 3797
rect -2854 3711 -2820 3729
rect -2854 3626 -2820 3661
rect -2596 5599 -2562 5634
rect -2596 5531 -2562 5549
rect -2596 5463 -2562 5477
rect -2596 5395 -2562 5405
rect -2596 5327 -2562 5333
rect -2596 5259 -2562 5261
rect -2596 5223 -2562 5225
rect -2596 5151 -2562 5157
rect -2596 5079 -2562 5089
rect -2596 5007 -2562 5021
rect -2596 4935 -2562 4953
rect -2596 4863 -2562 4885
rect -2596 4791 -2562 4817
rect -2596 4719 -2562 4749
rect -2596 4647 -2562 4681
rect -2596 4579 -2562 4613
rect -2596 4511 -2562 4541
rect -2596 4443 -2562 4469
rect -2596 4375 -2562 4397
rect -2596 4307 -2562 4325
rect -2596 4239 -2562 4253
rect -2596 4171 -2562 4181
rect -2596 4103 -2562 4109
rect -2596 4035 -2562 4037
rect -2596 3999 -2562 4001
rect -2596 3927 -2562 3933
rect -2596 3855 -2562 3865
rect -2596 3783 -2562 3797
rect -2596 3711 -2562 3729
rect -2596 3626 -2562 3661
rect -2154 5599 -2120 5634
rect -2154 5531 -2120 5549
rect -2154 5463 -2120 5477
rect -2154 5395 -2120 5405
rect -2154 5327 -2120 5333
rect -2154 5259 -2120 5261
rect -2154 5223 -2120 5225
rect -2154 5151 -2120 5157
rect -2154 5079 -2120 5089
rect -2154 5007 -2120 5021
rect -2154 4935 -2120 4953
rect -2154 4863 -2120 4885
rect -2154 4791 -2120 4817
rect -2154 4719 -2120 4749
rect -2154 4647 -2120 4681
rect -2154 4579 -2120 4613
rect -2154 4511 -2120 4541
rect -2154 4443 -2120 4469
rect -2154 4375 -2120 4397
rect -2154 4307 -2120 4325
rect -2154 4239 -2120 4253
rect -2154 4171 -2120 4181
rect -2154 4103 -2120 4109
rect -2154 4035 -2120 4037
rect -2154 3999 -2120 4001
rect -2154 3927 -2120 3933
rect -2154 3855 -2120 3865
rect -2154 3783 -2120 3797
rect -2154 3711 -2120 3729
rect -2154 3626 -2120 3661
rect -1896 5599 -1862 5634
rect -1896 5531 -1862 5549
rect -1896 5463 -1862 5477
rect -1896 5395 -1862 5405
rect -1896 5327 -1862 5333
rect -1896 5259 -1862 5261
rect -1896 5223 -1862 5225
rect -1896 5151 -1862 5157
rect -1896 5079 -1862 5089
rect -1896 5007 -1862 5021
rect -1896 4935 -1862 4953
rect -1896 4863 -1862 4885
rect -1896 4791 -1862 4817
rect -1896 4719 -1862 4749
rect -1896 4647 -1862 4681
rect -1896 4579 -1862 4613
rect -1896 4511 -1862 4541
rect -1896 4443 -1862 4469
rect -1896 4375 -1862 4397
rect -1896 4307 -1862 4325
rect -1896 4239 -1862 4253
rect -1896 4171 -1862 4181
rect -1896 4103 -1862 4109
rect -1896 4035 -1862 4037
rect -1896 3999 -1862 4001
rect -1896 3927 -1862 3933
rect -1896 3855 -1862 3865
rect -1896 3783 -1862 3797
rect -1896 3711 -1862 3729
rect -1896 3626 -1862 3661
rect -1454 5599 -1420 5634
rect -1454 5531 -1420 5549
rect -1454 5463 -1420 5477
rect -1454 5395 -1420 5405
rect -1454 5327 -1420 5333
rect -1454 5259 -1420 5261
rect -1454 5223 -1420 5225
rect -1454 5151 -1420 5157
rect -1454 5079 -1420 5089
rect -1454 5007 -1420 5021
rect -1454 4935 -1420 4953
rect -1454 4863 -1420 4885
rect -1454 4791 -1420 4817
rect -1454 4719 -1420 4749
rect -1454 4647 -1420 4681
rect -1454 4579 -1420 4613
rect -1454 4511 -1420 4541
rect -1454 4443 -1420 4469
rect -1454 4375 -1420 4397
rect -1454 4307 -1420 4325
rect -1454 4239 -1420 4253
rect -1454 4171 -1420 4181
rect -1454 4103 -1420 4109
rect -1454 4035 -1420 4037
rect -1454 3999 -1420 4001
rect -1454 3927 -1420 3933
rect -1454 3855 -1420 3865
rect -1454 3783 -1420 3797
rect -1454 3711 -1420 3729
rect -1454 3626 -1420 3661
rect -1196 5599 -1162 5634
rect -1196 5531 -1162 5549
rect -1196 5463 -1162 5477
rect -1196 5395 -1162 5405
rect -1196 5327 -1162 5333
rect -1196 5259 -1162 5261
rect -1196 5223 -1162 5225
rect -1196 5151 -1162 5157
rect -1196 5079 -1162 5089
rect -1196 5007 -1162 5021
rect -1196 4935 -1162 4953
rect -1196 4863 -1162 4885
rect -1196 4791 -1162 4817
rect -1196 4719 -1162 4749
rect -1196 4647 -1162 4681
rect -1196 4579 -1162 4613
rect -1196 4511 -1162 4541
rect -1196 4443 -1162 4469
rect -1196 4375 -1162 4397
rect -1196 4307 -1162 4325
rect -1196 4239 -1162 4253
rect -1196 4171 -1162 4181
rect -1196 4103 -1162 4109
rect -1196 4035 -1162 4037
rect -1196 3999 -1162 4001
rect -1196 3927 -1162 3933
rect -1196 3855 -1162 3865
rect -1196 3783 -1162 3797
rect -1196 3711 -1162 3729
rect -1196 3626 -1162 3661
rect -754 5599 -720 5634
rect -754 5531 -720 5549
rect -754 5463 -720 5477
rect -754 5395 -720 5405
rect -754 5327 -720 5333
rect -754 5259 -720 5261
rect -754 5223 -720 5225
rect -754 5151 -720 5157
rect -754 5079 -720 5089
rect -754 5007 -720 5021
rect -754 4935 -720 4953
rect -754 4863 -720 4885
rect -754 4791 -720 4817
rect -754 4719 -720 4749
rect -754 4647 -720 4681
rect -754 4579 -720 4613
rect -754 4511 -720 4541
rect -754 4443 -720 4469
rect -754 4375 -720 4397
rect -754 4307 -720 4325
rect -754 4239 -720 4253
rect -754 4171 -720 4181
rect -754 4103 -720 4109
rect -754 4035 -720 4037
rect -754 3999 -720 4001
rect -754 3927 -720 3933
rect -754 3855 -720 3865
rect -754 3783 -720 3797
rect -754 3711 -720 3729
rect -754 3626 -720 3661
rect -496 5599 -462 5634
rect -496 5531 -462 5549
rect -496 5463 -462 5477
rect -496 5395 -462 5405
rect -496 5327 -462 5333
rect -496 5259 -462 5261
rect -496 5223 -462 5225
rect -496 5151 -462 5157
rect -496 5079 -462 5089
rect -496 5007 -462 5021
rect -496 4935 -462 4953
rect -496 4863 -462 4885
rect -496 4791 -462 4817
rect -496 4719 -462 4749
rect -496 4647 -462 4681
rect -496 4579 -462 4613
rect -496 4511 -462 4541
rect -496 4443 -462 4469
rect -496 4375 -462 4397
rect -496 4307 -462 4325
rect -496 4239 -462 4253
rect -496 4171 -462 4181
rect -496 4103 -462 4109
rect -496 4035 -462 4037
rect -496 3999 -462 4001
rect -496 3927 -462 3933
rect -496 3855 -462 3865
rect -496 3783 -462 3797
rect -496 3711 -462 3729
rect -496 3626 -462 3661
rect -54 5599 -20 5634
rect -54 5531 -20 5549
rect -54 5463 -20 5477
rect -54 5395 -20 5405
rect -54 5327 -20 5333
rect -54 5259 -20 5261
rect -54 5223 -20 5225
rect -54 5151 -20 5157
rect -54 5079 -20 5089
rect -54 5007 -20 5021
rect -54 4935 -20 4953
rect -54 4863 -20 4885
rect -54 4791 -20 4817
rect -54 4719 -20 4749
rect -54 4647 -20 4681
rect -54 4579 -20 4613
rect -54 4511 -20 4541
rect -54 4443 -20 4469
rect -54 4375 -20 4397
rect -54 4307 -20 4325
rect -54 4239 -20 4253
rect -54 4171 -20 4181
rect -54 4103 -20 4109
rect -54 4035 -20 4037
rect -54 3999 -20 4001
rect -54 3927 -20 3933
rect -54 3855 -20 3865
rect -54 3783 -20 3797
rect -54 3711 -20 3729
rect -54 3626 -20 3661
rect 204 5599 238 5634
rect 204 5531 238 5549
rect 204 5463 238 5477
rect 204 5395 238 5405
rect 204 5327 238 5333
rect 204 5259 238 5261
rect 204 5223 238 5225
rect 204 5151 238 5157
rect 204 5079 238 5089
rect 204 5007 238 5021
rect 204 4935 238 4953
rect 204 4863 238 4885
rect 204 4791 238 4817
rect 204 4719 238 4749
rect 204 4647 238 4681
rect 204 4579 238 4613
rect 204 4511 238 4541
rect 204 4443 238 4469
rect 204 4375 238 4397
rect 204 4307 238 4325
rect 204 4239 238 4253
rect 204 4171 238 4181
rect 204 4103 238 4109
rect 204 4035 238 4037
rect 204 3999 238 4001
rect 204 3927 238 3933
rect 204 3855 238 3865
rect 204 3783 238 3797
rect 204 3711 238 3729
rect 204 3626 238 3661
rect 646 5599 680 5634
rect 646 5531 680 5549
rect 646 5463 680 5477
rect 646 5395 680 5405
rect 646 5327 680 5333
rect 646 5259 680 5261
rect 646 5223 680 5225
rect 646 5151 680 5157
rect 646 5079 680 5089
rect 646 5007 680 5021
rect 646 4935 680 4953
rect 646 4863 680 4885
rect 646 4791 680 4817
rect 646 4719 680 4749
rect 646 4647 680 4681
rect 646 4579 680 4613
rect 646 4511 680 4541
rect 646 4443 680 4469
rect 646 4375 680 4397
rect 646 4307 680 4325
rect 646 4239 680 4253
rect 646 4171 680 4181
rect 646 4103 680 4109
rect 646 4035 680 4037
rect 646 3999 680 4001
rect 646 3927 680 3933
rect 646 3855 680 3865
rect 646 3783 680 3797
rect 646 3711 680 3729
rect 646 3626 680 3661
rect 904 5599 938 5634
rect 904 5531 938 5549
rect 904 5463 938 5477
rect 904 5395 938 5405
rect 904 5327 938 5333
rect 904 5259 938 5261
rect 904 5223 938 5225
rect 904 5151 938 5157
rect 904 5079 938 5089
rect 904 5007 938 5021
rect 904 4935 938 4953
rect 904 4863 938 4885
rect 904 4791 938 4817
rect 904 4719 938 4749
rect 904 4647 938 4681
rect 904 4579 938 4613
rect 904 4511 938 4541
rect 904 4443 938 4469
rect 904 4375 938 4397
rect 904 4307 938 4325
rect 904 4239 938 4253
rect 904 4171 938 4181
rect 904 4103 938 4109
rect 904 4035 938 4037
rect 904 3999 938 4001
rect 904 3927 938 3933
rect 904 3855 938 3865
rect 904 3783 938 3797
rect 904 3711 938 3729
rect 904 3626 938 3661
rect 1346 5599 1380 5634
rect 1346 5531 1380 5549
rect 1346 5463 1380 5477
rect 1346 5395 1380 5405
rect 1346 5327 1380 5333
rect 1346 5259 1380 5261
rect 1346 5223 1380 5225
rect 1346 5151 1380 5157
rect 1346 5079 1380 5089
rect 1346 5007 1380 5021
rect 1346 4935 1380 4953
rect 1346 4863 1380 4885
rect 1346 4791 1380 4817
rect 1346 4719 1380 4749
rect 1346 4647 1380 4681
rect 1346 4579 1380 4613
rect 1346 4511 1380 4541
rect 1346 4443 1380 4469
rect 1346 4375 1380 4397
rect 1346 4307 1380 4325
rect 1346 4239 1380 4253
rect 1346 4171 1380 4181
rect 1346 4103 1380 4109
rect 1346 4035 1380 4037
rect 1346 3999 1380 4001
rect 1346 3927 1380 3933
rect 1346 3855 1380 3865
rect 1346 3783 1380 3797
rect 1346 3711 1380 3729
rect 1346 3626 1380 3661
rect 1604 5599 1638 5634
rect 1604 5531 1638 5549
rect 1604 5463 1638 5477
rect 1604 5395 1638 5405
rect 1604 5327 1638 5333
rect 1604 5259 1638 5261
rect 1604 5223 1638 5225
rect 1604 5151 1638 5157
rect 1604 5079 1638 5089
rect 1604 5007 1638 5021
rect 1604 4935 1638 4953
rect 1604 4863 1638 4885
rect 1604 4791 1638 4817
rect 1604 4719 1638 4749
rect 1604 4647 1638 4681
rect 1604 4579 1638 4613
rect 1604 4511 1638 4541
rect 1604 4443 1638 4469
rect 1604 4375 1638 4397
rect 1604 4307 1638 4325
rect 1604 4239 1638 4253
rect 1604 4171 1638 4181
rect 1604 4103 1638 4109
rect 1604 4035 1638 4037
rect 1604 3999 1638 4001
rect 1604 3927 1638 3933
rect 1604 3855 1638 3865
rect 1604 3783 1638 3797
rect 1604 3711 1638 3729
rect 1604 3626 1638 3661
rect 2046 5599 2080 5634
rect 2046 5531 2080 5549
rect 2046 5463 2080 5477
rect 2046 5395 2080 5405
rect 2046 5327 2080 5333
rect 2046 5259 2080 5261
rect 2046 5223 2080 5225
rect 2046 5151 2080 5157
rect 2046 5079 2080 5089
rect 2046 5007 2080 5021
rect 2046 4935 2080 4953
rect 2046 4863 2080 4885
rect 2046 4791 2080 4817
rect 2046 4719 2080 4749
rect 2046 4647 2080 4681
rect 2046 4579 2080 4613
rect 2046 4511 2080 4541
rect 2046 4443 2080 4469
rect 2046 4375 2080 4397
rect 2046 4307 2080 4325
rect 2046 4239 2080 4253
rect 2046 4171 2080 4181
rect 2046 4103 2080 4109
rect 2046 4035 2080 4037
rect 2046 3999 2080 4001
rect 2046 3927 2080 3933
rect 2046 3855 2080 3865
rect 2046 3783 2080 3797
rect 2046 3711 2080 3729
rect 2046 3626 2080 3661
rect 2304 5599 2338 5634
rect 2304 5531 2338 5549
rect 2304 5463 2338 5477
rect 2304 5395 2338 5405
rect 2304 5327 2338 5333
rect 2304 5259 2338 5261
rect 2304 5223 2338 5225
rect 2304 5151 2338 5157
rect 2304 5079 2338 5089
rect 2304 5007 2338 5021
rect 2304 4935 2338 4953
rect 2304 4863 2338 4885
rect 2304 4791 2338 4817
rect 2304 4719 2338 4749
rect 2304 4647 2338 4681
rect 2304 4579 2338 4613
rect 2304 4511 2338 4541
rect 2304 4443 2338 4469
rect 2304 4375 2338 4397
rect 2304 4307 2338 4325
rect 2304 4239 2338 4253
rect 2304 4171 2338 4181
rect 2304 4103 2338 4109
rect 2304 4035 2338 4037
rect 2304 3999 2338 4001
rect 2304 3927 2338 3933
rect 2304 3855 2338 3865
rect 2304 3783 2338 3797
rect 2304 3711 2338 3729
rect 2304 3626 2338 3661
rect 3746 5599 3780 5634
rect 3746 5531 3780 5549
rect 3746 5463 3780 5477
rect 3746 5395 3780 5405
rect 3746 5327 3780 5333
rect 3746 5259 3780 5261
rect 3746 5223 3780 5225
rect 3746 5151 3780 5157
rect 3746 5079 3780 5089
rect 3746 5007 3780 5021
rect 3746 4935 3780 4953
rect 3746 4863 3780 4885
rect 3746 4791 3780 4817
rect 3746 4719 3780 4749
rect 3746 4647 3780 4681
rect 3746 4579 3780 4613
rect 3746 4511 3780 4541
rect 3746 4443 3780 4469
rect 3746 4375 3780 4397
rect 3746 4307 3780 4325
rect 3746 4239 3780 4253
rect 3746 4171 3780 4181
rect 3746 4103 3780 4109
rect 3746 4035 3780 4037
rect 3746 3999 3780 4001
rect 3746 3927 3780 3933
rect 3746 3855 3780 3865
rect 3746 3783 3780 3797
rect 3746 3711 3780 3729
rect 3746 3626 3780 3661
rect 4004 5599 4038 5634
rect 4004 5531 4038 5549
rect 4004 5463 4038 5477
rect 4004 5395 4038 5405
rect 4004 5327 4038 5333
rect 4004 5259 4038 5261
rect 4004 5223 4038 5225
rect 4004 5151 4038 5157
rect 4004 5079 4038 5089
rect 4004 5007 4038 5021
rect 4004 4935 4038 4953
rect 4004 4863 4038 4885
rect 4004 4791 4038 4817
rect 4004 4719 4038 4749
rect 4004 4647 4038 4681
rect 4004 4579 4038 4613
rect 4004 4511 4038 4541
rect 4004 4443 4038 4469
rect 4004 4375 4038 4397
rect 4004 4307 4038 4325
rect 4004 4239 4038 4253
rect 4004 4171 4038 4181
rect 4004 4103 4038 4109
rect 4004 4035 4038 4037
rect 4004 3999 4038 4001
rect 4004 3927 4038 3933
rect 4004 3855 4038 3865
rect 4004 3783 4038 3797
rect 4004 3711 4038 3729
rect 4004 3626 4038 3661
rect 4446 5599 4480 5634
rect 4446 5531 4480 5549
rect 4446 5463 4480 5477
rect 4446 5395 4480 5405
rect 4446 5327 4480 5333
rect 4446 5259 4480 5261
rect 4446 5223 4480 5225
rect 4446 5151 4480 5157
rect 4446 5079 4480 5089
rect 4446 5007 4480 5021
rect 4446 4935 4480 4953
rect 4446 4863 4480 4885
rect 4446 4791 4480 4817
rect 4446 4719 4480 4749
rect 4446 4647 4480 4681
rect 4446 4579 4480 4613
rect 4446 4511 4480 4541
rect 4446 4443 4480 4469
rect 4446 4375 4480 4397
rect 4446 4307 4480 4325
rect 4446 4239 4480 4253
rect 4446 4171 4480 4181
rect 4446 4103 4480 4109
rect 4446 4035 4480 4037
rect 4446 3999 4480 4001
rect 4446 3927 4480 3933
rect 4446 3855 4480 3865
rect 4446 3783 4480 3797
rect 4446 3711 4480 3729
rect 4446 3626 4480 3661
rect 4704 5599 4738 5634
rect 4704 5531 4738 5549
rect 4704 5463 4738 5477
rect 4704 5395 4738 5405
rect 4704 5327 4738 5333
rect 4704 5259 4738 5261
rect 4704 5223 4738 5225
rect 4704 5151 4738 5157
rect 4704 5079 4738 5089
rect 4704 5007 4738 5021
rect 4704 4935 4738 4953
rect 4704 4863 4738 4885
rect 4704 4791 4738 4817
rect 4704 4719 4738 4749
rect 4704 4647 4738 4681
rect 4704 4579 4738 4613
rect 4704 4511 4738 4541
rect 4704 4443 4738 4469
rect 4704 4375 4738 4397
rect 4704 4307 4738 4325
rect 4704 4239 4738 4253
rect 4704 4171 4738 4181
rect 4704 4103 4738 4109
rect 4704 4035 4738 4037
rect 4704 3999 4738 4001
rect 4704 3927 4738 3933
rect 4704 3855 4738 3865
rect 4704 3783 4738 3797
rect 4704 3711 4738 3729
rect 4704 3626 4738 3661
rect 5146 5599 5180 5634
rect 5146 5531 5180 5549
rect 5146 5463 5180 5477
rect 5146 5395 5180 5405
rect 5146 5327 5180 5333
rect 5146 5259 5180 5261
rect 5146 5223 5180 5225
rect 5146 5151 5180 5157
rect 5146 5079 5180 5089
rect 5146 5007 5180 5021
rect 5146 4935 5180 4953
rect 5146 4863 5180 4885
rect 5146 4791 5180 4817
rect 5146 4719 5180 4749
rect 5146 4647 5180 4681
rect 5146 4579 5180 4613
rect 5146 4511 5180 4541
rect 5146 4443 5180 4469
rect 5146 4375 5180 4397
rect 5146 4307 5180 4325
rect 5146 4239 5180 4253
rect 5146 4171 5180 4181
rect 5146 4103 5180 4109
rect 5146 4035 5180 4037
rect 5146 3999 5180 4001
rect 5146 3927 5180 3933
rect 5146 3855 5180 3865
rect 5146 3783 5180 3797
rect 5146 3711 5180 3729
rect 5146 3626 5180 3661
rect 5404 5599 5438 5634
rect 5404 5531 5438 5549
rect 5404 5463 5438 5477
rect 5404 5395 5438 5405
rect 5404 5327 5438 5333
rect 5404 5259 5438 5261
rect 5404 5223 5438 5225
rect 5404 5151 5438 5157
rect 5404 5079 5438 5089
rect 5404 5007 5438 5021
rect 5404 4935 5438 4953
rect 5404 4863 5438 4885
rect 5404 4791 5438 4817
rect 5404 4719 5438 4749
rect 5404 4647 5438 4681
rect 5404 4579 5438 4613
rect 5404 4511 5438 4541
rect 5404 4443 5438 4469
rect 5404 4375 5438 4397
rect 5404 4307 5438 4325
rect 5404 4239 5438 4253
rect 5404 4171 5438 4181
rect 5404 4103 5438 4109
rect 5404 4035 5438 4037
rect 5404 3999 5438 4001
rect 5404 3927 5438 3933
rect 5404 3855 5438 3865
rect 5404 3783 5438 3797
rect 5404 3711 5438 3729
rect 5404 3626 5438 3661
rect 5846 5599 5880 5634
rect 5846 5531 5880 5549
rect 5846 5463 5880 5477
rect 5846 5395 5880 5405
rect 5846 5327 5880 5333
rect 5846 5259 5880 5261
rect 5846 5223 5880 5225
rect 5846 5151 5880 5157
rect 5846 5079 5880 5089
rect 5846 5007 5880 5021
rect 5846 4935 5880 4953
rect 5846 4863 5880 4885
rect 5846 4791 5880 4817
rect 5846 4719 5880 4749
rect 5846 4647 5880 4681
rect 5846 4579 5880 4613
rect 5846 4511 5880 4541
rect 5846 4443 5880 4469
rect 5846 4375 5880 4397
rect 5846 4307 5880 4325
rect 5846 4239 5880 4253
rect 5846 4171 5880 4181
rect 5846 4103 5880 4109
rect 5846 4035 5880 4037
rect 5846 3999 5880 4001
rect 5846 3927 5880 3933
rect 5846 3855 5880 3865
rect 5846 3783 5880 3797
rect 5846 3711 5880 3729
rect 5846 3626 5880 3661
rect 6104 5599 6138 5634
rect 6104 5531 6138 5549
rect 6104 5463 6138 5477
rect 6104 5395 6138 5405
rect 6104 5327 6138 5333
rect 6104 5259 6138 5261
rect 6104 5223 6138 5225
rect 6104 5151 6138 5157
rect 6104 5079 6138 5089
rect 6104 5007 6138 5021
rect 6104 4935 6138 4953
rect 6104 4863 6138 4885
rect 6104 4791 6138 4817
rect 6104 4719 6138 4749
rect 6104 4647 6138 4681
rect 6104 4579 6138 4613
rect 6104 4511 6138 4541
rect 6104 4443 6138 4469
rect 6104 4375 6138 4397
rect 6104 4307 6138 4325
rect 6104 4239 6138 4253
rect 6104 4171 6138 4181
rect 6104 4103 6138 4109
rect 6104 4035 6138 4037
rect 6104 3999 6138 4001
rect 6104 3927 6138 3933
rect 6104 3855 6138 3865
rect 6104 3783 6138 3797
rect 6104 3711 6138 3729
rect 6104 3626 6138 3661
rect 6546 5599 6580 5634
rect 6546 5531 6580 5549
rect 6546 5463 6580 5477
rect 6546 5395 6580 5405
rect 6546 5327 6580 5333
rect 6546 5259 6580 5261
rect 6546 5223 6580 5225
rect 6546 5151 6580 5157
rect 6546 5079 6580 5089
rect 6546 5007 6580 5021
rect 6546 4935 6580 4953
rect 6546 4863 6580 4885
rect 6546 4791 6580 4817
rect 6546 4719 6580 4749
rect 6546 4647 6580 4681
rect 6546 4579 6580 4613
rect 6546 4511 6580 4541
rect 6546 4443 6580 4469
rect 6546 4375 6580 4397
rect 6546 4307 6580 4325
rect 6546 4239 6580 4253
rect 6546 4171 6580 4181
rect 6546 4103 6580 4109
rect 6546 4035 6580 4037
rect 6546 3999 6580 4001
rect 6546 3927 6580 3933
rect 6546 3855 6580 3865
rect 6546 3783 6580 3797
rect 6546 3711 6580 3729
rect 6546 3626 6580 3661
rect 6804 5599 6838 5634
rect 6804 5531 6838 5549
rect 6804 5463 6838 5477
rect 6804 5395 6838 5405
rect 6804 5327 6838 5333
rect 6804 5259 6838 5261
rect 6804 5223 6838 5225
rect 6804 5151 6838 5157
rect 6804 5079 6838 5089
rect 6804 5007 6838 5021
rect 6804 4935 6838 4953
rect 6804 4863 6838 4885
rect 6804 4791 6838 4817
rect 6804 4719 6838 4749
rect 6804 4647 6838 4681
rect 6804 4579 6838 4613
rect 6804 4511 6838 4541
rect 6804 4443 6838 4469
rect 6804 4375 6838 4397
rect 6804 4307 6838 4325
rect 6804 4239 6838 4253
rect 6804 4171 6838 4181
rect 6804 4103 6838 4109
rect 6804 4035 6838 4037
rect 6804 3999 6838 4001
rect 6804 3927 6838 3933
rect 6804 3855 6838 3865
rect 6804 3783 6838 3797
rect 6804 3711 6838 3729
rect 6804 3626 6838 3661
rect 7246 5599 7280 5634
rect 7246 5531 7280 5549
rect 7246 5463 7280 5477
rect 7246 5395 7280 5405
rect 7246 5327 7280 5333
rect 7246 5259 7280 5261
rect 7246 5223 7280 5225
rect 7246 5151 7280 5157
rect 7246 5079 7280 5089
rect 7246 5007 7280 5021
rect 7246 4935 7280 4953
rect 7246 4863 7280 4885
rect 7246 4791 7280 4817
rect 7246 4719 7280 4749
rect 7246 4647 7280 4681
rect 7246 4579 7280 4613
rect 7246 4511 7280 4541
rect 7246 4443 7280 4469
rect 7246 4375 7280 4397
rect 7246 4307 7280 4325
rect 7246 4239 7280 4253
rect 7246 4171 7280 4181
rect 7246 4103 7280 4109
rect 7246 4035 7280 4037
rect 7246 3999 7280 4001
rect 7246 3927 7280 3933
rect 7246 3855 7280 3865
rect 7246 3783 7280 3797
rect 7246 3711 7280 3729
rect 7246 3626 7280 3661
rect 7504 5599 7538 5634
rect 7504 5531 7538 5549
rect 7504 5463 7538 5477
rect 7504 5395 7538 5405
rect 7504 5327 7538 5333
rect 7504 5259 7538 5261
rect 7504 5223 7538 5225
rect 7504 5151 7538 5157
rect 7504 5079 7538 5089
rect 7504 5007 7538 5021
rect 7504 4935 7538 4953
rect 7504 4863 7538 4885
rect 7504 4791 7538 4817
rect 7504 4719 7538 4749
rect 7504 4647 7538 4681
rect 7504 4579 7538 4613
rect 7504 4511 7538 4541
rect 7504 4443 7538 4469
rect 7504 4375 7538 4397
rect 7504 4307 7538 4325
rect 7504 4239 7538 4253
rect 7504 4171 7538 4181
rect 7504 4103 7538 4109
rect 7504 4035 7538 4037
rect 7504 3999 7538 4001
rect 7504 3927 7538 3933
rect 7504 3855 7538 3865
rect 7504 3783 7538 3797
rect 7504 3711 7538 3729
rect 7504 3626 7538 3661
rect 7946 5599 7980 5634
rect 7946 5531 7980 5549
rect 7946 5463 7980 5477
rect 7946 5395 7980 5405
rect 7946 5327 7980 5333
rect 7946 5259 7980 5261
rect 7946 5223 7980 5225
rect 7946 5151 7980 5157
rect 7946 5079 7980 5089
rect 7946 5007 7980 5021
rect 7946 4935 7980 4953
rect 7946 4863 7980 4885
rect 7946 4791 7980 4817
rect 7946 4719 7980 4749
rect 7946 4647 7980 4681
rect 7946 4579 7980 4613
rect 7946 4511 7980 4541
rect 7946 4443 7980 4469
rect 7946 4375 7980 4397
rect 7946 4307 7980 4325
rect 7946 4239 7980 4253
rect 7946 4171 7980 4181
rect 7946 4103 7980 4109
rect 7946 4035 7980 4037
rect 7946 3999 7980 4001
rect 7946 3927 7980 3933
rect 7946 3855 7980 3865
rect 7946 3783 7980 3797
rect 7946 3711 7980 3729
rect 7946 3626 7980 3661
rect 8204 5599 8238 5634
rect 8204 5531 8238 5549
rect 8204 5463 8238 5477
rect 8204 5395 8238 5405
rect 8204 5327 8238 5333
rect 8204 5259 8238 5261
rect 8204 5223 8238 5225
rect 8204 5151 8238 5157
rect 8204 5079 8238 5089
rect 8204 5007 8238 5021
rect 8204 4935 8238 4953
rect 8204 4863 8238 4885
rect 8204 4791 8238 4817
rect 8204 4719 8238 4749
rect 8204 4647 8238 4681
rect 8204 4579 8238 4613
rect 8204 4511 8238 4541
rect 8204 4443 8238 4469
rect 8204 4375 8238 4397
rect 8204 4307 8238 4325
rect 8204 4239 8238 4253
rect 8204 4171 8238 4181
rect 8204 4103 8238 4109
rect 8204 4035 8238 4037
rect 8204 3999 8238 4001
rect 8204 3927 8238 3933
rect 8204 3855 8238 3865
rect 8204 3783 8238 3797
rect 8204 3711 8238 3729
rect 8204 3626 8238 3661
rect 8646 5599 8680 5634
rect 8646 5531 8680 5549
rect 8646 5463 8680 5477
rect 8646 5395 8680 5405
rect 8646 5327 8680 5333
rect 8646 5259 8680 5261
rect 8646 5223 8680 5225
rect 8646 5151 8680 5157
rect 8646 5079 8680 5089
rect 8646 5007 8680 5021
rect 8646 4935 8680 4953
rect 8646 4863 8680 4885
rect 8646 4791 8680 4817
rect 8646 4719 8680 4749
rect 8646 4647 8680 4681
rect 8646 4579 8680 4613
rect 8646 4511 8680 4541
rect 8646 4443 8680 4469
rect 8646 4375 8680 4397
rect 8646 4307 8680 4325
rect 8646 4239 8680 4253
rect 8646 4171 8680 4181
rect 8646 4103 8680 4109
rect 8646 4035 8680 4037
rect 8646 3999 8680 4001
rect 8646 3927 8680 3933
rect 8646 3855 8680 3865
rect 8646 3783 8680 3797
rect 8646 3711 8680 3729
rect 8646 3626 8680 3661
rect 8904 5599 8938 5634
rect 8904 5531 8938 5549
rect 8904 5463 8938 5477
rect 8904 5395 8938 5405
rect 8904 5327 8938 5333
rect 8904 5259 8938 5261
rect 8904 5223 8938 5225
rect 8904 5151 8938 5157
rect 8904 5079 8938 5089
rect 8904 5007 8938 5021
rect 8904 4935 8938 4953
rect 8904 4863 8938 4885
rect 8904 4791 8938 4817
rect 8904 4719 8938 4749
rect 8904 4647 8938 4681
rect 8904 4579 8938 4613
rect 8904 4511 8938 4541
rect 8904 4443 8938 4469
rect 8904 4375 8938 4397
rect 8904 4307 8938 4325
rect 8904 4239 8938 4253
rect 8904 4171 8938 4181
rect 8904 4103 8938 4109
rect 8904 4035 8938 4037
rect 8904 3999 8938 4001
rect 8904 3927 8938 3933
rect 8904 3855 8938 3865
rect 8904 3783 8938 3797
rect 8904 3711 8938 3729
rect 8904 3626 8938 3661
rect 9346 5599 9380 5634
rect 9346 5531 9380 5549
rect 9346 5463 9380 5477
rect 9346 5395 9380 5405
rect 9346 5327 9380 5333
rect 9346 5259 9380 5261
rect 9346 5223 9380 5225
rect 9346 5151 9380 5157
rect 9346 5079 9380 5089
rect 9346 5007 9380 5021
rect 9346 4935 9380 4953
rect 9346 4863 9380 4885
rect 9346 4791 9380 4817
rect 9346 4719 9380 4749
rect 9346 4647 9380 4681
rect 9346 4579 9380 4613
rect 9346 4511 9380 4541
rect 9346 4443 9380 4469
rect 9346 4375 9380 4397
rect 9346 4307 9380 4325
rect 9346 4239 9380 4253
rect 9346 4171 9380 4181
rect 9346 4103 9380 4109
rect 9346 4035 9380 4037
rect 9346 3999 9380 4001
rect 9346 3927 9380 3933
rect 9346 3855 9380 3865
rect 9346 3783 9380 3797
rect 9346 3711 9380 3729
rect 9346 3626 9380 3661
rect 9604 5599 9638 5634
rect 9604 5531 9638 5549
rect 9604 5463 9638 5477
rect 9604 5395 9638 5405
rect 9604 5327 9638 5333
rect 9604 5259 9638 5261
rect 9604 5223 9638 5225
rect 9604 5151 9638 5157
rect 9604 5079 9638 5089
rect 9604 5007 9638 5021
rect 9604 4935 9638 4953
rect 9604 4863 9638 4885
rect 9604 4791 9638 4817
rect 9604 4719 9638 4749
rect 9604 4647 9638 4681
rect 9604 4579 9638 4613
rect 9604 4511 9638 4541
rect 9604 4443 9638 4469
rect 9604 4375 9638 4397
rect 9604 4307 9638 4325
rect 9604 4239 9638 4253
rect 9604 4171 9638 4181
rect 9604 4103 9638 4109
rect 9604 4035 9638 4037
rect 9604 3999 9638 4001
rect 9604 3927 9638 3933
rect 9604 3855 9638 3865
rect 9604 3783 9638 3797
rect 9604 3711 9638 3729
rect 9604 3626 9638 3661
rect 10046 5599 10080 5634
rect 10046 5531 10080 5549
rect 10046 5463 10080 5477
rect 10046 5395 10080 5405
rect 10046 5327 10080 5333
rect 10046 5259 10080 5261
rect 10046 5223 10080 5225
rect 10046 5151 10080 5157
rect 10046 5079 10080 5089
rect 10046 5007 10080 5021
rect 10046 4935 10080 4953
rect 10046 4863 10080 4885
rect 10046 4791 10080 4817
rect 10046 4719 10080 4749
rect 10046 4647 10080 4681
rect 10046 4579 10080 4613
rect 10046 4511 10080 4541
rect 10046 4443 10080 4469
rect 10046 4375 10080 4397
rect 10046 4307 10080 4325
rect 10046 4239 10080 4253
rect 10046 4171 10080 4181
rect 10046 4103 10080 4109
rect 10046 4035 10080 4037
rect 10046 3999 10080 4001
rect 10046 3927 10080 3933
rect 10046 3855 10080 3865
rect 10046 3783 10080 3797
rect 10046 3711 10080 3729
rect 10046 3626 10080 3661
rect 10304 5599 10338 5634
rect 11742 5628 11781 5662
rect 11823 5628 11853 5662
rect 11891 5628 11925 5662
rect 11959 5628 11993 5662
rect 12031 5628 12061 5662
rect 12103 5628 12142 5662
rect 12642 5628 12681 5662
rect 12723 5628 12753 5662
rect 12791 5628 12825 5662
rect 12859 5628 12893 5662
rect 12931 5628 12961 5662
rect 13003 5628 13042 5662
rect 13542 5628 13581 5662
rect 13623 5628 13653 5662
rect 13691 5628 13725 5662
rect 13759 5628 13793 5662
rect 13831 5628 13861 5662
rect 13903 5628 13942 5662
rect 14442 5628 14481 5662
rect 14523 5628 14553 5662
rect 14591 5628 14625 5662
rect 14659 5628 14693 5662
rect 14731 5628 14761 5662
rect 14803 5628 14842 5662
rect 15342 5628 15381 5662
rect 15423 5628 15453 5662
rect 15491 5628 15525 5662
rect 15559 5628 15593 5662
rect 15631 5628 15661 5662
rect 15703 5628 15742 5662
rect 16242 5628 16281 5662
rect 16323 5628 16353 5662
rect 16391 5628 16425 5662
rect 16459 5628 16493 5662
rect 16531 5628 16561 5662
rect 16603 5628 16642 5662
rect 17142 5628 17181 5662
rect 17223 5628 17253 5662
rect 17291 5628 17325 5662
rect 17359 5628 17393 5662
rect 17431 5628 17461 5662
rect 17503 5628 17542 5662
rect 18042 5628 18081 5662
rect 18123 5628 18153 5662
rect 18191 5628 18225 5662
rect 18259 5628 18293 5662
rect 18331 5628 18361 5662
rect 18403 5628 18442 5662
rect 10304 5531 10338 5549
rect 10304 5463 10338 5477
rect 11866 5489 12004 5505
rect 11866 5455 11882 5489
rect 11916 5455 11954 5489
rect 11988 5455 12004 5489
rect 11866 5439 12004 5455
rect 12766 5489 12904 5505
rect 12766 5455 12782 5489
rect 12816 5455 12854 5489
rect 12888 5455 12904 5489
rect 12766 5439 12904 5455
rect 13666 5489 13804 5505
rect 13666 5455 13682 5489
rect 13716 5455 13754 5489
rect 13788 5455 13804 5489
rect 13666 5439 13804 5455
rect 14566 5489 14704 5505
rect 14566 5455 14582 5489
rect 14616 5455 14654 5489
rect 14688 5455 14704 5489
rect 14566 5439 14704 5455
rect 15466 5489 15604 5505
rect 15466 5455 15482 5489
rect 15516 5455 15554 5489
rect 15588 5455 15604 5489
rect 15466 5439 15604 5455
rect 16366 5489 16504 5505
rect 16366 5455 16382 5489
rect 16416 5455 16454 5489
rect 16488 5455 16504 5489
rect 16366 5439 16504 5455
rect 17266 5489 17404 5505
rect 17266 5455 17282 5489
rect 17316 5455 17354 5489
rect 17388 5455 17404 5489
rect 17266 5439 17404 5455
rect 18166 5489 18304 5505
rect 18166 5455 18182 5489
rect 18216 5455 18254 5489
rect 18288 5455 18304 5489
rect 18166 5439 18304 5455
rect 10304 5395 10338 5405
rect 10304 5327 10338 5333
rect 10304 5259 10338 5261
rect 10304 5223 10338 5225
rect 10304 5151 10338 5157
rect 10304 5079 10338 5089
rect 10304 5007 10338 5021
rect 10304 4935 10338 4953
rect 10304 4863 10338 4885
rect 10304 4791 10338 4817
rect 10304 4719 10338 4749
rect 10304 4647 10338 4681
rect 10304 4579 10338 4613
rect 10304 4511 10338 4541
rect 10304 4443 10338 4469
rect 10304 4375 10338 4397
rect 10304 4307 10338 4325
rect 10304 4239 10338 4253
rect 10304 4171 10338 4181
rect 10304 4103 10338 4109
rect 10304 4035 10338 4037
rect 10304 3999 10338 4001
rect 10304 3927 10338 3933
rect 10304 3855 10338 3865
rect 10304 3783 10338 3797
rect 10304 3711 10338 3729
rect 10304 3626 10338 3661
rect -4208 3558 -4161 3592
rect -4125 3558 -4091 3592
rect -4055 3558 -4008 3592
rect -3508 3558 -3461 3592
rect -3425 3558 -3391 3592
rect -3355 3558 -3308 3592
rect -2808 3558 -2761 3592
rect -2725 3558 -2691 3592
rect -2655 3558 -2608 3592
rect -2108 3558 -2061 3592
rect -2025 3558 -1991 3592
rect -1955 3558 -1908 3592
rect -1408 3558 -1361 3592
rect -1325 3558 -1291 3592
rect -1255 3558 -1208 3592
rect -708 3558 -661 3592
rect -625 3558 -591 3592
rect -555 3558 -508 3592
rect -8 3558 39 3592
rect 75 3558 109 3592
rect 145 3558 192 3592
rect 692 3558 739 3592
rect 775 3558 809 3592
rect 845 3558 892 3592
rect 1392 3558 1439 3592
rect 1475 3558 1509 3592
rect 1545 3558 1592 3592
rect 2092 3558 2139 3592
rect 2175 3558 2209 3592
rect 2245 3558 2292 3592
rect 3792 3558 3839 3592
rect 3875 3558 3909 3592
rect 3945 3558 3992 3592
rect 4492 3558 4539 3592
rect 4575 3558 4609 3592
rect 4645 3558 4692 3592
rect 5192 3558 5239 3592
rect 5275 3558 5309 3592
rect 5345 3558 5392 3592
rect 5892 3558 5939 3592
rect 5975 3558 6009 3592
rect 6045 3558 6092 3592
rect 6592 3558 6639 3592
rect 6675 3558 6709 3592
rect 6745 3558 6792 3592
rect 7292 3558 7339 3592
rect 7375 3558 7409 3592
rect 7445 3558 7492 3592
rect 7992 3558 8039 3592
rect 8075 3558 8109 3592
rect 8145 3558 8192 3592
rect 8692 3558 8739 3592
rect 8775 3558 8809 3592
rect 8845 3558 8892 3592
rect 9392 3558 9439 3592
rect 9475 3558 9509 3592
rect 9545 3558 9592 3592
rect 10092 3558 10139 3592
rect 10175 3558 10209 3592
rect 10245 3558 10292 3592
rect 1269 2134 1407 2150
rect 1269 2100 1285 2134
rect 1319 2100 1357 2134
rect 1391 2100 1407 2134
rect 1269 2084 1407 2100
rect 2269 2134 2407 2150
rect 2269 2100 2285 2134
rect 2319 2100 2357 2134
rect 2391 2100 2407 2134
rect 2269 2084 2407 2100
rect 3269 2134 3407 2150
rect 3269 2100 3285 2134
rect 3319 2100 3357 2134
rect 3391 2100 3407 2134
rect 3269 2084 3407 2100
rect 4269 2134 4407 2150
rect 4269 2100 4285 2134
rect 4319 2100 4357 2134
rect 4391 2100 4407 2134
rect 4269 2084 4407 2100
rect 5269 2134 5407 2150
rect 5269 2100 5285 2134
rect 5319 2100 5357 2134
rect 5391 2100 5407 2134
rect 5269 2084 5407 2100
rect 6269 2134 6407 2150
rect 6269 2100 6285 2134
rect 6319 2100 6357 2134
rect 6391 2100 6407 2134
rect 6269 2084 6407 2100
rect 7269 2134 7407 2150
rect 7269 2100 7285 2134
rect 7319 2100 7357 2134
rect 7391 2100 7407 2134
rect 7269 2084 7407 2100
rect 8269 2134 8407 2150
rect 8269 2100 8285 2134
rect 8319 2100 8357 2134
rect 8391 2100 8407 2134
rect 8269 2084 8407 2100
rect 9269 2134 9407 2150
rect 9269 2100 9285 2134
rect 9319 2100 9357 2134
rect 9391 2100 9407 2134
rect 9269 2084 9407 2100
rect 10269 2134 10407 2150
rect 10269 2100 10285 2134
rect 10319 2100 10357 2134
rect 10391 2100 10407 2134
rect 10269 2084 10407 2100
rect 1134 1954 1173 1988
rect 1215 1954 1245 1988
rect 1283 1954 1317 1988
rect 1351 1954 1385 1988
rect 1423 1954 1453 1988
rect 1495 1954 1534 1988
rect 2134 1954 2173 1988
rect 2215 1954 2245 1988
rect 2283 1954 2317 1988
rect 2351 1954 2385 1988
rect 2423 1954 2453 1988
rect 2495 1954 2534 1988
rect 3134 1954 3173 1988
rect 3215 1954 3245 1988
rect 3283 1954 3317 1988
rect 3351 1954 3385 1988
rect 3423 1954 3453 1988
rect 3495 1954 3534 1988
rect 4134 1954 4173 1988
rect 4215 1954 4245 1988
rect 4283 1954 4317 1988
rect 4351 1954 4385 1988
rect 4423 1954 4453 1988
rect 4495 1954 4534 1988
rect 5134 1954 5173 1988
rect 5215 1954 5245 1988
rect 5283 1954 5317 1988
rect 5351 1954 5385 1988
rect 5423 1954 5453 1988
rect 5495 1954 5534 1988
rect 6134 1954 6173 1988
rect 6215 1954 6245 1988
rect 6283 1954 6317 1988
rect 6351 1954 6385 1988
rect 6423 1954 6453 1988
rect 6495 1954 6534 1988
rect 7134 1954 7173 1988
rect 7215 1954 7245 1988
rect 7283 1954 7317 1988
rect 7351 1954 7385 1988
rect 7423 1954 7453 1988
rect 7495 1954 7534 1988
rect 8134 1954 8173 1988
rect 8215 1954 8245 1988
rect 8283 1954 8317 1988
rect 8351 1954 8385 1988
rect 8423 1954 8453 1988
rect 8495 1954 8534 1988
rect 9134 1954 9173 1988
rect 9215 1954 9245 1988
rect 9283 1954 9317 1988
rect 9351 1954 9385 1988
rect 9423 1954 9453 1988
rect 9495 1954 9534 1988
rect 10134 1954 10173 1988
rect 10215 1954 10245 1988
rect 10283 1954 10317 1988
rect 10351 1954 10385 1988
rect 10423 1954 10453 1988
rect 10495 1954 10534 1988
rect 1088 1901 1122 1920
rect 1088 1833 1122 1835
rect 1088 1797 1122 1799
rect 1088 1712 1122 1731
rect 1546 1901 1580 1920
rect 1546 1833 1580 1835
rect 1546 1797 1580 1799
rect 1546 1712 1580 1731
rect 2088 1901 2122 1920
rect 2088 1833 2122 1835
rect 2088 1797 2122 1799
rect 2088 1712 2122 1731
rect 2546 1901 2580 1920
rect 2546 1833 2580 1835
rect 2546 1797 2580 1799
rect 2546 1712 2580 1731
rect 3088 1901 3122 1920
rect 3088 1833 3122 1835
rect 3088 1797 3122 1799
rect 3088 1712 3122 1731
rect 3546 1901 3580 1920
rect 3546 1833 3580 1835
rect 3546 1797 3580 1799
rect 3546 1712 3580 1731
rect 4088 1901 4122 1920
rect 4088 1833 4122 1835
rect 4088 1797 4122 1799
rect 4088 1712 4122 1731
rect 4546 1901 4580 1920
rect 4546 1833 4580 1835
rect 4546 1797 4580 1799
rect 4546 1712 4580 1731
rect 5088 1901 5122 1920
rect 5088 1833 5122 1835
rect 5088 1797 5122 1799
rect 5088 1712 5122 1731
rect 5546 1901 5580 1920
rect 5546 1833 5580 1835
rect 5546 1797 5580 1799
rect 5546 1712 5580 1731
rect 6088 1901 6122 1920
rect 6088 1833 6122 1835
rect 6088 1797 6122 1799
rect 6088 1712 6122 1731
rect 6546 1901 6580 1920
rect 6546 1833 6580 1835
rect 6546 1797 6580 1799
rect 6546 1712 6580 1731
rect 7088 1901 7122 1920
rect 7088 1833 7122 1835
rect 7088 1797 7122 1799
rect 7088 1712 7122 1731
rect 7546 1901 7580 1920
rect 7546 1833 7580 1835
rect 7546 1797 7580 1799
rect 7546 1712 7580 1731
rect 8088 1901 8122 1920
rect 8088 1833 8122 1835
rect 8088 1797 8122 1799
rect 8088 1712 8122 1731
rect 8546 1901 8580 1920
rect 8546 1833 8580 1835
rect 8546 1797 8580 1799
rect 8546 1712 8580 1731
rect 9088 1901 9122 1920
rect 9088 1833 9122 1835
rect 9088 1797 9122 1799
rect 9088 1712 9122 1731
rect 9546 1901 9580 1920
rect 9546 1833 9580 1835
rect 9546 1797 9580 1799
rect 9546 1712 9580 1731
rect 10088 1901 10122 1920
rect 10088 1833 10122 1835
rect 10088 1797 10122 1799
rect 10088 1712 10122 1731
rect 10546 1901 10580 1920
rect 10546 1833 10580 1835
rect 10546 1797 10580 1799
rect 10546 1712 10580 1731
rect 1134 1644 1173 1678
rect 1215 1644 1245 1678
rect 1283 1644 1317 1678
rect 1351 1644 1385 1678
rect 1423 1644 1453 1678
rect 1495 1644 1534 1678
rect 2134 1644 2173 1678
rect 2215 1644 2245 1678
rect 2283 1644 2317 1678
rect 2351 1644 2385 1678
rect 2423 1644 2453 1678
rect 2495 1644 2534 1678
rect 3134 1644 3173 1678
rect 3215 1644 3245 1678
rect 3283 1644 3317 1678
rect 3351 1644 3385 1678
rect 3423 1644 3453 1678
rect 3495 1644 3534 1678
rect 4134 1644 4173 1678
rect 4215 1644 4245 1678
rect 4283 1644 4317 1678
rect 4351 1644 4385 1678
rect 4423 1644 4453 1678
rect 4495 1644 4534 1678
rect 5134 1644 5173 1678
rect 5215 1644 5245 1678
rect 5283 1644 5317 1678
rect 5351 1644 5385 1678
rect 5423 1644 5453 1678
rect 5495 1644 5534 1678
rect 6134 1644 6173 1678
rect 6215 1644 6245 1678
rect 6283 1644 6317 1678
rect 6351 1644 6385 1678
rect 6423 1644 6453 1678
rect 6495 1644 6534 1678
rect 7134 1644 7173 1678
rect 7215 1644 7245 1678
rect 7283 1644 7317 1678
rect 7351 1644 7385 1678
rect 7423 1644 7453 1678
rect 7495 1644 7534 1678
rect 8134 1644 8173 1678
rect 8215 1644 8245 1678
rect 8283 1644 8317 1678
rect 8351 1644 8385 1678
rect 8423 1644 8453 1678
rect 8495 1644 8534 1678
rect 9134 1644 9173 1678
rect 9215 1644 9245 1678
rect 9283 1644 9317 1678
rect 9351 1644 9385 1678
rect 9423 1644 9453 1678
rect 9495 1644 9534 1678
rect 10134 1644 10173 1678
rect 10215 1644 10245 1678
rect 10283 1644 10317 1678
rect 10351 1644 10385 1678
rect 10423 1644 10453 1678
rect 10495 1644 10534 1678
rect 1134 1454 1173 1488
rect 1215 1454 1245 1488
rect 1283 1454 1317 1488
rect 1351 1454 1385 1488
rect 1423 1454 1453 1488
rect 1495 1454 1534 1488
rect 2134 1454 2173 1488
rect 2215 1454 2245 1488
rect 2283 1454 2317 1488
rect 2351 1454 2385 1488
rect 2423 1454 2453 1488
rect 2495 1454 2534 1488
rect 3134 1454 3173 1488
rect 3215 1454 3245 1488
rect 3283 1454 3317 1488
rect 3351 1454 3385 1488
rect 3423 1454 3453 1488
rect 3495 1454 3534 1488
rect 4134 1454 4173 1488
rect 4215 1454 4245 1488
rect 4283 1454 4317 1488
rect 4351 1454 4385 1488
rect 4423 1454 4453 1488
rect 4495 1454 4534 1488
rect 5134 1454 5173 1488
rect 5215 1454 5245 1488
rect 5283 1454 5317 1488
rect 5351 1454 5385 1488
rect 5423 1454 5453 1488
rect 5495 1454 5534 1488
rect 6134 1454 6173 1488
rect 6215 1454 6245 1488
rect 6283 1454 6317 1488
rect 6351 1454 6385 1488
rect 6423 1454 6453 1488
rect 6495 1454 6534 1488
rect 7134 1454 7173 1488
rect 7215 1454 7245 1488
rect 7283 1454 7317 1488
rect 7351 1454 7385 1488
rect 7423 1454 7453 1488
rect 7495 1454 7534 1488
rect 8134 1454 8173 1488
rect 8215 1454 8245 1488
rect 8283 1454 8317 1488
rect 8351 1454 8385 1488
rect 8423 1454 8453 1488
rect 8495 1454 8534 1488
rect 9134 1454 9173 1488
rect 9215 1454 9245 1488
rect 9283 1454 9317 1488
rect 9351 1454 9385 1488
rect 9423 1454 9453 1488
rect 9495 1454 9534 1488
rect 10134 1454 10173 1488
rect 10215 1454 10245 1488
rect 10283 1454 10317 1488
rect 10351 1454 10385 1488
rect 10423 1454 10453 1488
rect 10495 1454 10534 1488
rect 1088 1401 1122 1420
rect 1088 1333 1122 1335
rect 1088 1297 1122 1299
rect 1088 1212 1122 1231
rect 1546 1401 1580 1420
rect 1546 1333 1580 1335
rect 1546 1297 1580 1299
rect 1546 1212 1580 1231
rect 2088 1401 2122 1420
rect 2088 1333 2122 1335
rect 2088 1297 2122 1299
rect 2088 1212 2122 1231
rect 2546 1401 2580 1420
rect 2546 1333 2580 1335
rect 2546 1297 2580 1299
rect 2546 1212 2580 1231
rect 3088 1401 3122 1420
rect 3088 1333 3122 1335
rect 3088 1297 3122 1299
rect 3088 1212 3122 1231
rect 3546 1401 3580 1420
rect 3546 1333 3580 1335
rect 3546 1297 3580 1299
rect 3546 1212 3580 1231
rect 4088 1401 4122 1420
rect 4088 1333 4122 1335
rect 4088 1297 4122 1299
rect 4088 1212 4122 1231
rect 4546 1401 4580 1420
rect 4546 1333 4580 1335
rect 4546 1297 4580 1299
rect 4546 1212 4580 1231
rect 5088 1401 5122 1420
rect 5088 1333 5122 1335
rect 5088 1297 5122 1299
rect 5088 1212 5122 1231
rect 5546 1401 5580 1420
rect 5546 1333 5580 1335
rect 5546 1297 5580 1299
rect 5546 1212 5580 1231
rect 6088 1401 6122 1420
rect 6088 1333 6122 1335
rect 6088 1297 6122 1299
rect 6088 1212 6122 1231
rect 6546 1401 6580 1420
rect 6546 1333 6580 1335
rect 6546 1297 6580 1299
rect 6546 1212 6580 1231
rect 7088 1401 7122 1420
rect 7088 1333 7122 1335
rect 7088 1297 7122 1299
rect 7088 1212 7122 1231
rect 7546 1401 7580 1420
rect 7546 1333 7580 1335
rect 7546 1297 7580 1299
rect 7546 1212 7580 1231
rect 8088 1401 8122 1420
rect 8088 1333 8122 1335
rect 8088 1297 8122 1299
rect 8088 1212 8122 1231
rect 8546 1401 8580 1420
rect 8546 1333 8580 1335
rect 8546 1297 8580 1299
rect 8546 1212 8580 1231
rect 9088 1401 9122 1420
rect 9088 1333 9122 1335
rect 9088 1297 9122 1299
rect 9088 1212 9122 1231
rect 9546 1401 9580 1420
rect 9546 1333 9580 1335
rect 9546 1297 9580 1299
rect 9546 1212 9580 1231
rect 10088 1401 10122 1420
rect 10088 1333 10122 1335
rect 10088 1297 10122 1299
rect 10088 1212 10122 1231
rect 10546 1401 10580 1420
rect 10546 1333 10580 1335
rect 10546 1297 10580 1299
rect 10546 1212 10580 1231
rect 1134 1144 1173 1178
rect 1215 1144 1245 1178
rect 1283 1144 1317 1178
rect 1351 1144 1385 1178
rect 1423 1144 1453 1178
rect 1495 1144 1534 1178
rect 2134 1144 2173 1178
rect 2215 1144 2245 1178
rect 2283 1144 2317 1178
rect 2351 1144 2385 1178
rect 2423 1144 2453 1178
rect 2495 1144 2534 1178
rect 3134 1144 3173 1178
rect 3215 1144 3245 1178
rect 3283 1144 3317 1178
rect 3351 1144 3385 1178
rect 3423 1144 3453 1178
rect 3495 1144 3534 1178
rect 4134 1144 4173 1178
rect 4215 1144 4245 1178
rect 4283 1144 4317 1178
rect 4351 1144 4385 1178
rect 4423 1144 4453 1178
rect 4495 1144 4534 1178
rect 5134 1144 5173 1178
rect 5215 1144 5245 1178
rect 5283 1144 5317 1178
rect 5351 1144 5385 1178
rect 5423 1144 5453 1178
rect 5495 1144 5534 1178
rect 6134 1144 6173 1178
rect 6215 1144 6245 1178
rect 6283 1144 6317 1178
rect 6351 1144 6385 1178
rect 6423 1144 6453 1178
rect 6495 1144 6534 1178
rect 7134 1144 7173 1178
rect 7215 1144 7245 1178
rect 7283 1144 7317 1178
rect 7351 1144 7385 1178
rect 7423 1144 7453 1178
rect 7495 1144 7534 1178
rect 8134 1144 8173 1178
rect 8215 1144 8245 1178
rect 8283 1144 8317 1178
rect 8351 1144 8385 1178
rect 8423 1144 8453 1178
rect 8495 1144 8534 1178
rect 9134 1144 9173 1178
rect 9215 1144 9245 1178
rect 9283 1144 9317 1178
rect 9351 1144 9385 1178
rect 9423 1144 9453 1178
rect 9495 1144 9534 1178
rect 10134 1144 10173 1178
rect 10215 1144 10245 1178
rect 10283 1144 10317 1178
rect 10351 1144 10385 1178
rect 10423 1144 10453 1178
rect 10495 1144 10534 1178
rect 1268 997 1406 1013
rect 1268 963 1284 997
rect 1318 963 1356 997
rect 1390 963 1406 997
rect 1268 947 1406 963
rect 2268 997 2406 1013
rect 2268 963 2284 997
rect 2318 963 2356 997
rect 2390 963 2406 997
rect 2268 947 2406 963
rect 3268 997 3406 1013
rect 3268 963 3284 997
rect 3318 963 3356 997
rect 3390 963 3406 997
rect 3268 947 3406 963
rect 4268 997 4406 1013
rect 4268 963 4284 997
rect 4318 963 4356 997
rect 4390 963 4406 997
rect 4268 947 4406 963
rect 5268 997 5406 1013
rect 5268 963 5284 997
rect 5318 963 5356 997
rect 5390 963 5406 997
rect 5268 947 5406 963
rect 6268 997 6406 1013
rect 6268 963 6284 997
rect 6318 963 6356 997
rect 6390 963 6406 997
rect 6268 947 6406 963
rect 7268 997 7406 1013
rect 7268 963 7284 997
rect 7318 963 7356 997
rect 7390 963 7406 997
rect 7268 947 7406 963
rect 8268 997 8406 1013
rect 8268 963 8284 997
rect 8318 963 8356 997
rect 8390 963 8406 997
rect 8268 947 8406 963
rect 9268 997 9406 1013
rect 9268 963 9284 997
rect 9318 963 9356 997
rect 9390 963 9406 997
rect 9268 947 9406 963
rect 10268 997 10406 1013
rect 10268 963 10284 997
rect 10318 963 10356 997
rect 10390 963 10406 997
rect 10268 947 10406 963
<< viali >>
rect 2167 8720 2201 8754
rect 2239 8720 2273 8754
rect 3167 8720 3201 8754
rect 3239 8720 3273 8754
rect 2063 8556 2071 8590
rect 2071 8556 2097 8590
rect 2135 8556 2139 8590
rect 2139 8556 2169 8590
rect 2207 8556 2241 8590
rect 2279 8556 2309 8590
rect 2309 8556 2313 8590
rect 2351 8556 2377 8590
rect 2377 8556 2385 8590
rect 3063 8556 3071 8590
rect 3071 8556 3097 8590
rect 3135 8556 3139 8590
rect 3139 8556 3169 8590
rect 3207 8556 3241 8590
rect 3279 8556 3309 8590
rect 3309 8556 3313 8590
rect 3351 8556 3377 8590
rect 3377 8556 3385 8590
rect 1978 8462 2012 8470
rect 1978 8436 2012 8462
rect 1978 8394 2012 8398
rect 1978 8364 2012 8394
rect 1978 8292 2012 8326
rect 1978 8224 2012 8254
rect 1978 8220 2012 8224
rect 1978 8156 2012 8182
rect 1978 8148 2012 8156
rect 2436 8462 2470 8470
rect 2436 8436 2470 8462
rect 2436 8394 2470 8398
rect 2436 8364 2470 8394
rect 2436 8292 2470 8326
rect 2436 8224 2470 8254
rect 2436 8220 2470 8224
rect 2436 8156 2470 8182
rect 2436 8148 2470 8156
rect 2978 8462 3012 8470
rect 2978 8436 3012 8462
rect 2978 8394 3012 8398
rect 2978 8364 3012 8394
rect 2978 8292 3012 8326
rect 2978 8224 3012 8254
rect 2978 8220 3012 8224
rect 2978 8156 3012 8182
rect 2978 8148 3012 8156
rect 21455 8506 21561 8900
rect 3436 8462 3470 8470
rect 3436 8436 3470 8462
rect 3436 8394 3470 8398
rect 3436 8364 3470 8394
rect 3436 8292 3470 8326
rect 3436 8224 3470 8254
rect 3436 8220 3470 8224
rect 3436 8156 3470 8182
rect 3436 8148 3470 8156
rect 2063 8028 2071 8062
rect 2071 8028 2097 8062
rect 2135 8028 2139 8062
rect 2139 8028 2169 8062
rect 2207 8028 2241 8062
rect 2279 8028 2309 8062
rect 2309 8028 2313 8062
rect 2351 8028 2377 8062
rect 2377 8028 2385 8062
rect 3063 8028 3071 8062
rect 3071 8028 3097 8062
rect 3135 8028 3139 8062
rect 3139 8028 3169 8062
rect 3207 8028 3241 8062
rect 3279 8028 3309 8062
rect 3309 8028 3313 8062
rect 3351 8028 3377 8062
rect 3377 8028 3385 8062
rect 2063 7816 2071 7850
rect 2071 7816 2097 7850
rect 2135 7816 2139 7850
rect 2139 7816 2169 7850
rect 2207 7816 2241 7850
rect 2279 7816 2309 7850
rect 2309 7816 2313 7850
rect 2351 7816 2377 7850
rect 2377 7816 2385 7850
rect 3063 7816 3071 7850
rect 3071 7816 3097 7850
rect 3135 7816 3139 7850
rect 3139 7816 3169 7850
rect 3207 7816 3241 7850
rect 3279 7816 3309 7850
rect 3309 7816 3313 7850
rect 3351 7816 3377 7850
rect 3377 7816 3385 7850
rect 1978 7722 2012 7730
rect 1978 7696 2012 7722
rect 1978 7654 2012 7658
rect 1978 7624 2012 7654
rect 1978 7552 2012 7586
rect 1978 7484 2012 7514
rect 1978 7480 2012 7484
rect 1978 7416 2012 7442
rect 1978 7408 2012 7416
rect 2436 7722 2470 7730
rect 2436 7696 2470 7722
rect 2436 7654 2470 7658
rect 2436 7624 2470 7654
rect 2436 7552 2470 7586
rect 2436 7484 2470 7514
rect 2436 7480 2470 7484
rect 2436 7416 2470 7442
rect 2436 7408 2470 7416
rect 2978 7722 3012 7730
rect 2978 7696 3012 7722
rect 2978 7654 3012 7658
rect 2978 7624 3012 7654
rect 2978 7552 3012 7586
rect 2978 7484 3012 7514
rect 2978 7480 3012 7484
rect 2978 7416 3012 7442
rect 2978 7408 3012 7416
rect 3436 7722 3470 7730
rect 3436 7696 3470 7722
rect 3436 7654 3470 7658
rect 3436 7624 3470 7654
rect 3436 7552 3470 7586
rect 3436 7484 3470 7514
rect 3436 7480 3470 7484
rect 21097 7569 21131 7602
rect 21097 7568 21131 7569
rect 21097 7497 21131 7530
rect 21097 7496 21131 7497
rect 3436 7416 3470 7442
rect 3436 7408 3470 7416
rect 2063 7288 2071 7322
rect 2071 7288 2097 7322
rect 2135 7288 2139 7322
rect 2139 7288 2169 7322
rect 2207 7288 2241 7322
rect 2279 7288 2309 7322
rect 2309 7288 2313 7322
rect 2351 7288 2377 7322
rect 2377 7288 2385 7322
rect 3063 7288 3071 7322
rect 3071 7288 3097 7322
rect 3135 7288 3139 7322
rect 3139 7288 3169 7322
rect 3207 7288 3241 7322
rect 3279 7288 3309 7322
rect 3309 7288 3313 7322
rect 3351 7288 3377 7322
rect 3377 7288 3385 7322
rect 2164 7115 2198 7149
rect 2236 7115 2270 7149
rect 3164 7115 3198 7149
rect 3236 7115 3270 7149
rect 11885 7060 11919 7094
rect 11957 7060 11991 7094
rect 12785 7060 12819 7094
rect 12857 7060 12891 7094
rect 13685 7060 13719 7094
rect 13757 7060 13791 7094
rect 14585 7060 14619 7094
rect 14657 7060 14691 7094
rect 15485 7060 15519 7094
rect 15557 7060 15591 7094
rect 16385 7060 16419 7094
rect 16457 7060 16491 7094
rect 17285 7060 17319 7094
rect 17357 7060 17391 7094
rect 18185 7060 18219 7094
rect 18257 7060 18291 7094
rect 11781 6896 11789 6930
rect 11789 6896 11815 6930
rect 11853 6896 11857 6930
rect 11857 6896 11887 6930
rect 11925 6896 11959 6930
rect 11997 6896 12027 6930
rect 12027 6896 12031 6930
rect 12069 6896 12095 6930
rect 12095 6896 12103 6930
rect 12681 6896 12689 6930
rect 12689 6896 12715 6930
rect 12753 6896 12757 6930
rect 12757 6896 12787 6930
rect 12825 6896 12859 6930
rect 12897 6896 12927 6930
rect 12927 6896 12931 6930
rect 12969 6896 12995 6930
rect 12995 6896 13003 6930
rect 13581 6896 13589 6930
rect 13589 6896 13615 6930
rect 13653 6896 13657 6930
rect 13657 6896 13687 6930
rect 13725 6896 13759 6930
rect 13797 6896 13827 6930
rect 13827 6896 13831 6930
rect 13869 6896 13895 6930
rect 13895 6896 13903 6930
rect 14481 6896 14489 6930
rect 14489 6896 14515 6930
rect 14553 6896 14557 6930
rect 14557 6896 14587 6930
rect 14625 6896 14659 6930
rect 14697 6896 14727 6930
rect 14727 6896 14731 6930
rect 14769 6896 14795 6930
rect 14795 6896 14803 6930
rect 15381 6896 15389 6930
rect 15389 6896 15415 6930
rect 15453 6896 15457 6930
rect 15457 6896 15487 6930
rect 15525 6896 15559 6930
rect 15597 6896 15627 6930
rect 15627 6896 15631 6930
rect 15669 6896 15695 6930
rect 15695 6896 15703 6930
rect 16281 6896 16289 6930
rect 16289 6896 16315 6930
rect 16353 6896 16357 6930
rect 16357 6896 16387 6930
rect 16425 6896 16459 6930
rect 16497 6896 16527 6930
rect 16527 6896 16531 6930
rect 16569 6896 16595 6930
rect 16595 6896 16603 6930
rect 17181 6896 17189 6930
rect 17189 6896 17215 6930
rect 17253 6896 17257 6930
rect 17257 6896 17287 6930
rect 17325 6896 17359 6930
rect 17397 6896 17427 6930
rect 17427 6896 17431 6930
rect 17469 6896 17495 6930
rect 17495 6896 17503 6930
rect 18081 6896 18089 6930
rect 18089 6896 18115 6930
rect 18153 6896 18157 6930
rect 18157 6896 18187 6930
rect 18225 6896 18259 6930
rect 18297 6896 18327 6930
rect 18327 6896 18331 6930
rect 18369 6896 18395 6930
rect 18395 6896 18403 6930
rect 11696 6802 11730 6810
rect 11696 6776 11730 6802
rect 11696 6734 11730 6738
rect 11696 6704 11730 6734
rect 11696 6632 11730 6666
rect 11696 6564 11730 6594
rect 11696 6560 11730 6564
rect 11696 6496 11730 6522
rect 11696 6488 11730 6496
rect 12154 6802 12188 6810
rect 12154 6776 12188 6802
rect 12154 6734 12188 6738
rect 12154 6704 12188 6734
rect 12154 6632 12188 6666
rect 12154 6564 12188 6594
rect 12154 6560 12188 6564
rect 12154 6496 12188 6522
rect 12154 6488 12188 6496
rect 12596 6802 12630 6810
rect 12596 6776 12630 6802
rect 12596 6734 12630 6738
rect 12596 6704 12630 6734
rect 12596 6632 12630 6666
rect 12596 6564 12630 6594
rect 12596 6560 12630 6564
rect 12596 6496 12630 6522
rect 12596 6488 12630 6496
rect 13054 6802 13088 6810
rect 13054 6776 13088 6802
rect 13054 6734 13088 6738
rect 13054 6704 13088 6734
rect 13054 6632 13088 6666
rect 13054 6564 13088 6594
rect 13054 6560 13088 6564
rect 13054 6496 13088 6522
rect 13054 6488 13088 6496
rect 13496 6802 13530 6810
rect 13496 6776 13530 6802
rect 13496 6734 13530 6738
rect 13496 6704 13530 6734
rect 13496 6632 13530 6666
rect 13496 6564 13530 6594
rect 13496 6560 13530 6564
rect 13496 6496 13530 6522
rect 13496 6488 13530 6496
rect 13954 6802 13988 6810
rect 13954 6776 13988 6802
rect 13954 6734 13988 6738
rect 13954 6704 13988 6734
rect 13954 6632 13988 6666
rect 13954 6564 13988 6594
rect 13954 6560 13988 6564
rect 13954 6496 13988 6522
rect 13954 6488 13988 6496
rect 14396 6802 14430 6810
rect 14396 6776 14430 6802
rect 14396 6734 14430 6738
rect 14396 6704 14430 6734
rect 14396 6632 14430 6666
rect 14396 6564 14430 6594
rect 14396 6560 14430 6564
rect 14396 6496 14430 6522
rect 14396 6488 14430 6496
rect 14854 6802 14888 6810
rect 14854 6776 14888 6802
rect 14854 6734 14888 6738
rect 14854 6704 14888 6734
rect 14854 6632 14888 6666
rect 14854 6564 14888 6594
rect 14854 6560 14888 6564
rect 14854 6496 14888 6522
rect 14854 6488 14888 6496
rect 15296 6802 15330 6810
rect 15296 6776 15330 6802
rect 15296 6734 15330 6738
rect 15296 6704 15330 6734
rect 15296 6632 15330 6666
rect 15296 6564 15330 6594
rect 15296 6560 15330 6564
rect 15296 6496 15330 6522
rect 15296 6488 15330 6496
rect 15754 6802 15788 6810
rect 15754 6776 15788 6802
rect 15754 6734 15788 6738
rect 15754 6704 15788 6734
rect 15754 6632 15788 6666
rect 15754 6564 15788 6594
rect 15754 6560 15788 6564
rect 15754 6496 15788 6522
rect 15754 6488 15788 6496
rect 16196 6802 16230 6810
rect 16196 6776 16230 6802
rect 16196 6734 16230 6738
rect 16196 6704 16230 6734
rect 16196 6632 16230 6666
rect 16196 6564 16230 6594
rect 16196 6560 16230 6564
rect 16196 6496 16230 6522
rect 16196 6488 16230 6496
rect 16654 6802 16688 6810
rect 16654 6776 16688 6802
rect 16654 6734 16688 6738
rect 16654 6704 16688 6734
rect 16654 6632 16688 6666
rect 16654 6564 16688 6594
rect 16654 6560 16688 6564
rect 16654 6496 16688 6522
rect 16654 6488 16688 6496
rect 17096 6802 17130 6810
rect 17096 6776 17130 6802
rect 17096 6734 17130 6738
rect 17096 6704 17130 6734
rect 17096 6632 17130 6666
rect 17096 6564 17130 6594
rect 17096 6560 17130 6564
rect 17096 6496 17130 6522
rect 17096 6488 17130 6496
rect 17554 6802 17588 6810
rect 17554 6776 17588 6802
rect 17554 6734 17588 6738
rect 17554 6704 17588 6734
rect 17554 6632 17588 6666
rect 17554 6564 17588 6594
rect 17554 6560 17588 6564
rect 17554 6496 17588 6522
rect 17554 6488 17588 6496
rect 17996 6802 18030 6810
rect 17996 6776 18030 6802
rect 17996 6734 18030 6738
rect 17996 6704 18030 6734
rect 17996 6632 18030 6666
rect 17996 6564 18030 6594
rect 17996 6560 18030 6564
rect 17996 6496 18030 6522
rect 17996 6488 18030 6496
rect 18454 6802 18488 6810
rect 18454 6776 18488 6802
rect 18454 6734 18488 6738
rect 18454 6704 18488 6734
rect 18454 6632 18488 6666
rect 18454 6564 18488 6594
rect 18454 6560 18488 6564
rect 18454 6496 18488 6522
rect 18454 6488 18488 6496
rect 11781 6368 11789 6402
rect 11789 6368 11815 6402
rect 11853 6368 11857 6402
rect 11857 6368 11887 6402
rect 11925 6368 11959 6402
rect 11997 6368 12027 6402
rect 12027 6368 12031 6402
rect 12069 6368 12095 6402
rect 12095 6368 12103 6402
rect 12681 6368 12689 6402
rect 12689 6368 12715 6402
rect 12753 6368 12757 6402
rect 12757 6368 12787 6402
rect 12825 6368 12859 6402
rect 12897 6368 12927 6402
rect 12927 6368 12931 6402
rect 12969 6368 12995 6402
rect 12995 6368 13003 6402
rect 13581 6368 13589 6402
rect 13589 6368 13615 6402
rect 13653 6368 13657 6402
rect 13657 6368 13687 6402
rect 13725 6368 13759 6402
rect 13797 6368 13827 6402
rect 13827 6368 13831 6402
rect 13869 6368 13895 6402
rect 13895 6368 13903 6402
rect 14481 6368 14489 6402
rect 14489 6368 14515 6402
rect 14553 6368 14557 6402
rect 14557 6368 14587 6402
rect 14625 6368 14659 6402
rect 14697 6368 14727 6402
rect 14727 6368 14731 6402
rect 14769 6368 14795 6402
rect 14795 6368 14803 6402
rect 15381 6368 15389 6402
rect 15389 6368 15415 6402
rect 15453 6368 15457 6402
rect 15457 6368 15487 6402
rect 15525 6368 15559 6402
rect 15597 6368 15627 6402
rect 15627 6368 15631 6402
rect 15669 6368 15695 6402
rect 15695 6368 15703 6402
rect 16281 6368 16289 6402
rect 16289 6368 16315 6402
rect 16353 6368 16357 6402
rect 16357 6368 16387 6402
rect 16425 6368 16459 6402
rect 16497 6368 16527 6402
rect 16527 6368 16531 6402
rect 16569 6368 16595 6402
rect 16595 6368 16603 6402
rect 17181 6368 17189 6402
rect 17189 6368 17215 6402
rect 17253 6368 17257 6402
rect 17257 6368 17287 6402
rect 17325 6368 17359 6402
rect 17397 6368 17427 6402
rect 17427 6368 17431 6402
rect 17469 6368 17495 6402
rect 17495 6368 17503 6402
rect 18081 6368 18089 6402
rect 18089 6368 18115 6402
rect 18153 6368 18157 6402
rect 18157 6368 18187 6402
rect 18225 6368 18259 6402
rect 18297 6368 18327 6402
rect 18327 6368 18331 6402
rect 18369 6368 18395 6402
rect 18395 6368 18403 6402
rect 11781 6156 11789 6190
rect 11789 6156 11815 6190
rect 11853 6156 11857 6190
rect 11857 6156 11887 6190
rect 11925 6156 11959 6190
rect 11997 6156 12027 6190
rect 12027 6156 12031 6190
rect 12069 6156 12095 6190
rect 12095 6156 12103 6190
rect 12681 6156 12689 6190
rect 12689 6156 12715 6190
rect 12753 6156 12757 6190
rect 12757 6156 12787 6190
rect 12825 6156 12859 6190
rect 12897 6156 12927 6190
rect 12927 6156 12931 6190
rect 12969 6156 12995 6190
rect 12995 6156 13003 6190
rect 13581 6156 13589 6190
rect 13589 6156 13615 6190
rect 13653 6156 13657 6190
rect 13657 6156 13687 6190
rect 13725 6156 13759 6190
rect 13797 6156 13827 6190
rect 13827 6156 13831 6190
rect 13869 6156 13895 6190
rect 13895 6156 13903 6190
rect 14481 6156 14489 6190
rect 14489 6156 14515 6190
rect 14553 6156 14557 6190
rect 14557 6156 14587 6190
rect 14625 6156 14659 6190
rect 14697 6156 14727 6190
rect 14727 6156 14731 6190
rect 14769 6156 14795 6190
rect 14795 6156 14803 6190
rect 15381 6156 15389 6190
rect 15389 6156 15415 6190
rect 15453 6156 15457 6190
rect 15457 6156 15487 6190
rect 15525 6156 15559 6190
rect 15597 6156 15627 6190
rect 15627 6156 15631 6190
rect 15669 6156 15695 6190
rect 15695 6156 15703 6190
rect 16281 6156 16289 6190
rect 16289 6156 16315 6190
rect 16353 6156 16357 6190
rect 16357 6156 16387 6190
rect 16425 6156 16459 6190
rect 16497 6156 16527 6190
rect 16527 6156 16531 6190
rect 16569 6156 16595 6190
rect 16595 6156 16603 6190
rect 17181 6156 17189 6190
rect 17189 6156 17215 6190
rect 17253 6156 17257 6190
rect 17257 6156 17287 6190
rect 17325 6156 17359 6190
rect 17397 6156 17427 6190
rect 17427 6156 17431 6190
rect 17469 6156 17495 6190
rect 17495 6156 17503 6190
rect 18081 6156 18089 6190
rect 18089 6156 18115 6190
rect 18153 6156 18157 6190
rect 18157 6156 18187 6190
rect 18225 6156 18259 6190
rect 18297 6156 18327 6190
rect 18327 6156 18331 6190
rect 18369 6156 18395 6190
rect 18395 6156 18403 6190
rect 11696 6062 11730 6070
rect 11696 6036 11730 6062
rect 11696 5994 11730 5998
rect 11696 5964 11730 5994
rect 11696 5892 11730 5926
rect 11696 5824 11730 5854
rect 11696 5820 11730 5824
rect 11696 5756 11730 5782
rect 11696 5748 11730 5756
rect 12154 6062 12188 6070
rect 12154 6036 12188 6062
rect 12154 5994 12188 5998
rect 12154 5964 12188 5994
rect 12154 5892 12188 5926
rect 12154 5824 12188 5854
rect 12154 5820 12188 5824
rect 12154 5756 12188 5782
rect 12154 5748 12188 5756
rect 12596 6062 12630 6070
rect 12596 6036 12630 6062
rect 12596 5994 12630 5998
rect 12596 5964 12630 5994
rect 12596 5892 12630 5926
rect 12596 5824 12630 5854
rect 12596 5820 12630 5824
rect 12596 5756 12630 5782
rect 12596 5748 12630 5756
rect 13054 6062 13088 6070
rect 13054 6036 13088 6062
rect 13054 5994 13088 5998
rect 13054 5964 13088 5994
rect 13054 5892 13088 5926
rect 13054 5824 13088 5854
rect 13054 5820 13088 5824
rect 13054 5756 13088 5782
rect 13054 5748 13088 5756
rect 13496 6062 13530 6070
rect 13496 6036 13530 6062
rect 13496 5994 13530 5998
rect 13496 5964 13530 5994
rect 13496 5892 13530 5926
rect 13496 5824 13530 5854
rect 13496 5820 13530 5824
rect 13496 5756 13530 5782
rect 13496 5748 13530 5756
rect 13954 6062 13988 6070
rect 13954 6036 13988 6062
rect 13954 5994 13988 5998
rect 13954 5964 13988 5994
rect 13954 5892 13988 5926
rect 13954 5824 13988 5854
rect 13954 5820 13988 5824
rect 13954 5756 13988 5782
rect 13954 5748 13988 5756
rect 14396 6062 14430 6070
rect 14396 6036 14430 6062
rect 14396 5994 14430 5998
rect 14396 5964 14430 5994
rect 14396 5892 14430 5926
rect 14396 5824 14430 5854
rect 14396 5820 14430 5824
rect 14396 5756 14430 5782
rect 14396 5748 14430 5756
rect 14854 6062 14888 6070
rect 14854 6036 14888 6062
rect 14854 5994 14888 5998
rect 14854 5964 14888 5994
rect 14854 5892 14888 5926
rect 14854 5824 14888 5854
rect 14854 5820 14888 5824
rect 14854 5756 14888 5782
rect 14854 5748 14888 5756
rect 15296 6062 15330 6070
rect 15296 6036 15330 6062
rect 15296 5994 15330 5998
rect 15296 5964 15330 5994
rect 15296 5892 15330 5926
rect 15296 5824 15330 5854
rect 15296 5820 15330 5824
rect 15296 5756 15330 5782
rect 15296 5748 15330 5756
rect 15754 6062 15788 6070
rect 15754 6036 15788 6062
rect 15754 5994 15788 5998
rect 15754 5964 15788 5994
rect 15754 5892 15788 5926
rect 15754 5824 15788 5854
rect 15754 5820 15788 5824
rect 15754 5756 15788 5782
rect 15754 5748 15788 5756
rect 16196 6062 16230 6070
rect 16196 6036 16230 6062
rect 16196 5994 16230 5998
rect 16196 5964 16230 5994
rect 16196 5892 16230 5926
rect 16196 5824 16230 5854
rect 16196 5820 16230 5824
rect 16196 5756 16230 5782
rect 16196 5748 16230 5756
rect 16654 6062 16688 6070
rect 16654 6036 16688 6062
rect 16654 5994 16688 5998
rect 16654 5964 16688 5994
rect 16654 5892 16688 5926
rect 16654 5824 16688 5854
rect 16654 5820 16688 5824
rect 16654 5756 16688 5782
rect 16654 5748 16688 5756
rect 17096 6062 17130 6070
rect 17096 6036 17130 6062
rect 17096 5994 17130 5998
rect 17096 5964 17130 5994
rect 17096 5892 17130 5926
rect 17096 5824 17130 5854
rect 17096 5820 17130 5824
rect 17096 5756 17130 5782
rect 17096 5748 17130 5756
rect 17554 6062 17588 6070
rect 17554 6036 17588 6062
rect 17554 5994 17588 5998
rect 17554 5964 17588 5994
rect 17554 5892 17588 5926
rect 17554 5824 17588 5854
rect 17554 5820 17588 5824
rect 17554 5756 17588 5782
rect 17554 5748 17588 5756
rect 17996 6062 18030 6070
rect 17996 6036 18030 6062
rect 17996 5994 18030 5998
rect 17996 5964 18030 5994
rect 17996 5892 18030 5926
rect 17996 5824 18030 5854
rect 17996 5820 18030 5824
rect 17996 5756 18030 5782
rect 17996 5748 18030 5756
rect 18454 6062 18488 6070
rect 18454 6036 18488 6062
rect 21455 6075 21561 6469
rect 18454 5994 18488 5998
rect 18454 5964 18488 5994
rect 18454 5892 18488 5926
rect 18454 5824 18488 5854
rect 18454 5820 18488 5824
rect 18454 5756 18488 5782
rect 18454 5748 18488 5756
rect -4161 5668 -4159 5702
rect -4159 5668 -4127 5702
rect -4089 5668 -4057 5702
rect -4057 5668 -4055 5702
rect -3461 5668 -3459 5702
rect -3459 5668 -3427 5702
rect -3389 5668 -3357 5702
rect -3357 5668 -3355 5702
rect -2761 5668 -2759 5702
rect -2759 5668 -2727 5702
rect -2689 5668 -2657 5702
rect -2657 5668 -2655 5702
rect -2061 5668 -2059 5702
rect -2059 5668 -2027 5702
rect -1989 5668 -1957 5702
rect -1957 5668 -1955 5702
rect -1361 5668 -1359 5702
rect -1359 5668 -1327 5702
rect -1289 5668 -1257 5702
rect -1257 5668 -1255 5702
rect -661 5668 -659 5702
rect -659 5668 -627 5702
rect -589 5668 -557 5702
rect -557 5668 -555 5702
rect 39 5668 41 5702
rect 41 5668 73 5702
rect 111 5668 143 5702
rect 143 5668 145 5702
rect 739 5668 741 5702
rect 741 5668 773 5702
rect 811 5668 843 5702
rect 843 5668 845 5702
rect 1439 5668 1441 5702
rect 1441 5668 1473 5702
rect 1511 5668 1543 5702
rect 1543 5668 1545 5702
rect 2139 5668 2141 5702
rect 2141 5668 2173 5702
rect 2211 5668 2243 5702
rect 2243 5668 2245 5702
rect 3839 5668 3841 5702
rect 3841 5668 3873 5702
rect 3911 5668 3943 5702
rect 3943 5668 3945 5702
rect 4539 5668 4541 5702
rect 4541 5668 4573 5702
rect 4611 5668 4643 5702
rect 4643 5668 4645 5702
rect 5239 5668 5241 5702
rect 5241 5668 5273 5702
rect 5311 5668 5343 5702
rect 5343 5668 5345 5702
rect 5939 5668 5941 5702
rect 5941 5668 5973 5702
rect 6011 5668 6043 5702
rect 6043 5668 6045 5702
rect 6639 5668 6641 5702
rect 6641 5668 6673 5702
rect 6711 5668 6743 5702
rect 6743 5668 6745 5702
rect 7339 5668 7341 5702
rect 7341 5668 7373 5702
rect 7411 5668 7443 5702
rect 7443 5668 7445 5702
rect 8039 5668 8041 5702
rect 8041 5668 8073 5702
rect 8111 5668 8143 5702
rect 8143 5668 8145 5702
rect 8739 5668 8741 5702
rect 8741 5668 8773 5702
rect 8811 5668 8843 5702
rect 8843 5668 8845 5702
rect 9439 5668 9441 5702
rect 9441 5668 9473 5702
rect 9511 5668 9543 5702
rect 9543 5668 9545 5702
rect 10139 5668 10141 5702
rect 10141 5668 10173 5702
rect 10211 5668 10243 5702
rect 10243 5668 10245 5702
rect -4254 5565 -4220 5583
rect -4254 5549 -4220 5565
rect -4254 5497 -4220 5511
rect -4254 5477 -4220 5497
rect -4254 5429 -4220 5439
rect -4254 5405 -4220 5429
rect -4254 5361 -4220 5367
rect -4254 5333 -4220 5361
rect -4254 5293 -4220 5295
rect -4254 5261 -4220 5293
rect -4254 5191 -4220 5223
rect -4254 5189 -4220 5191
rect -4254 5123 -4220 5151
rect -4254 5117 -4220 5123
rect -4254 5055 -4220 5079
rect -4254 5045 -4220 5055
rect -4254 4987 -4220 5007
rect -4254 4973 -4220 4987
rect -4254 4919 -4220 4935
rect -4254 4901 -4220 4919
rect -4254 4851 -4220 4863
rect -4254 4829 -4220 4851
rect -4254 4783 -4220 4791
rect -4254 4757 -4220 4783
rect -4254 4715 -4220 4719
rect -4254 4685 -4220 4715
rect -4254 4613 -4220 4647
rect -4254 4545 -4220 4575
rect -4254 4541 -4220 4545
rect -4254 4477 -4220 4503
rect -4254 4469 -4220 4477
rect -4254 4409 -4220 4431
rect -4254 4397 -4220 4409
rect -4254 4341 -4220 4359
rect -4254 4325 -4220 4341
rect -4254 4273 -4220 4287
rect -4254 4253 -4220 4273
rect -4254 4205 -4220 4215
rect -4254 4181 -4220 4205
rect -4254 4137 -4220 4143
rect -4254 4109 -4220 4137
rect -4254 4069 -4220 4071
rect -4254 4037 -4220 4069
rect -4254 3967 -4220 3999
rect -4254 3965 -4220 3967
rect -4254 3899 -4220 3927
rect -4254 3893 -4220 3899
rect -4254 3831 -4220 3855
rect -4254 3821 -4220 3831
rect -4254 3763 -4220 3783
rect -4254 3749 -4220 3763
rect -4254 3695 -4220 3711
rect -4254 3677 -4220 3695
rect -3996 5565 -3962 5583
rect -3996 5549 -3962 5565
rect -3996 5497 -3962 5511
rect -3996 5477 -3962 5497
rect -3996 5429 -3962 5439
rect -3996 5405 -3962 5429
rect -3996 5361 -3962 5367
rect -3996 5333 -3962 5361
rect -3996 5293 -3962 5295
rect -3996 5261 -3962 5293
rect -3996 5191 -3962 5223
rect -3996 5189 -3962 5191
rect -3996 5123 -3962 5151
rect -3996 5117 -3962 5123
rect -3996 5055 -3962 5079
rect -3996 5045 -3962 5055
rect -3996 4987 -3962 5007
rect -3996 4973 -3962 4987
rect -3996 4919 -3962 4935
rect -3996 4901 -3962 4919
rect -3996 4851 -3962 4863
rect -3996 4829 -3962 4851
rect -3996 4783 -3962 4791
rect -3996 4757 -3962 4783
rect -3996 4715 -3962 4719
rect -3996 4685 -3962 4715
rect -3996 4613 -3962 4647
rect -3996 4545 -3962 4575
rect -3996 4541 -3962 4545
rect -3996 4477 -3962 4503
rect -3996 4469 -3962 4477
rect -3996 4409 -3962 4431
rect -3996 4397 -3962 4409
rect -3996 4341 -3962 4359
rect -3996 4325 -3962 4341
rect -3996 4273 -3962 4287
rect -3996 4253 -3962 4273
rect -3996 4205 -3962 4215
rect -3996 4181 -3962 4205
rect -3996 4137 -3962 4143
rect -3996 4109 -3962 4137
rect -3996 4069 -3962 4071
rect -3996 4037 -3962 4069
rect -3996 3967 -3962 3999
rect -3996 3965 -3962 3967
rect -3996 3899 -3962 3927
rect -3996 3893 -3962 3899
rect -3996 3831 -3962 3855
rect -3996 3821 -3962 3831
rect -3996 3763 -3962 3783
rect -3996 3749 -3962 3763
rect -3996 3695 -3962 3711
rect -3996 3677 -3962 3695
rect -3554 5565 -3520 5583
rect -3554 5549 -3520 5565
rect -3554 5497 -3520 5511
rect -3554 5477 -3520 5497
rect -3554 5429 -3520 5439
rect -3554 5405 -3520 5429
rect -3554 5361 -3520 5367
rect -3554 5333 -3520 5361
rect -3554 5293 -3520 5295
rect -3554 5261 -3520 5293
rect -3554 5191 -3520 5223
rect -3554 5189 -3520 5191
rect -3554 5123 -3520 5151
rect -3554 5117 -3520 5123
rect -3554 5055 -3520 5079
rect -3554 5045 -3520 5055
rect -3554 4987 -3520 5007
rect -3554 4973 -3520 4987
rect -3554 4919 -3520 4935
rect -3554 4901 -3520 4919
rect -3554 4851 -3520 4863
rect -3554 4829 -3520 4851
rect -3554 4783 -3520 4791
rect -3554 4757 -3520 4783
rect -3554 4715 -3520 4719
rect -3554 4685 -3520 4715
rect -3554 4613 -3520 4647
rect -3554 4545 -3520 4575
rect -3554 4541 -3520 4545
rect -3554 4477 -3520 4503
rect -3554 4469 -3520 4477
rect -3554 4409 -3520 4431
rect -3554 4397 -3520 4409
rect -3554 4341 -3520 4359
rect -3554 4325 -3520 4341
rect -3554 4273 -3520 4287
rect -3554 4253 -3520 4273
rect -3554 4205 -3520 4215
rect -3554 4181 -3520 4205
rect -3554 4137 -3520 4143
rect -3554 4109 -3520 4137
rect -3554 4069 -3520 4071
rect -3554 4037 -3520 4069
rect -3554 3967 -3520 3999
rect -3554 3965 -3520 3967
rect -3554 3899 -3520 3927
rect -3554 3893 -3520 3899
rect -3554 3831 -3520 3855
rect -3554 3821 -3520 3831
rect -3554 3763 -3520 3783
rect -3554 3749 -3520 3763
rect -3554 3695 -3520 3711
rect -3554 3677 -3520 3695
rect -3296 5565 -3262 5583
rect -3296 5549 -3262 5565
rect -3296 5497 -3262 5511
rect -3296 5477 -3262 5497
rect -3296 5429 -3262 5439
rect -3296 5405 -3262 5429
rect -3296 5361 -3262 5367
rect -3296 5333 -3262 5361
rect -3296 5293 -3262 5295
rect -3296 5261 -3262 5293
rect -3296 5191 -3262 5223
rect -3296 5189 -3262 5191
rect -3296 5123 -3262 5151
rect -3296 5117 -3262 5123
rect -3296 5055 -3262 5079
rect -3296 5045 -3262 5055
rect -3296 4987 -3262 5007
rect -3296 4973 -3262 4987
rect -3296 4919 -3262 4935
rect -3296 4901 -3262 4919
rect -3296 4851 -3262 4863
rect -3296 4829 -3262 4851
rect -3296 4783 -3262 4791
rect -3296 4757 -3262 4783
rect -3296 4715 -3262 4719
rect -3296 4685 -3262 4715
rect -3296 4613 -3262 4647
rect -3296 4545 -3262 4575
rect -3296 4541 -3262 4545
rect -3296 4477 -3262 4503
rect -3296 4469 -3262 4477
rect -3296 4409 -3262 4431
rect -3296 4397 -3262 4409
rect -3296 4341 -3262 4359
rect -3296 4325 -3262 4341
rect -3296 4273 -3262 4287
rect -3296 4253 -3262 4273
rect -3296 4205 -3262 4215
rect -3296 4181 -3262 4205
rect -3296 4137 -3262 4143
rect -3296 4109 -3262 4137
rect -3296 4069 -3262 4071
rect -3296 4037 -3262 4069
rect -3296 3967 -3262 3999
rect -3296 3965 -3262 3967
rect -3296 3899 -3262 3927
rect -3296 3893 -3262 3899
rect -3296 3831 -3262 3855
rect -3296 3821 -3262 3831
rect -3296 3763 -3262 3783
rect -3296 3749 -3262 3763
rect -3296 3695 -3262 3711
rect -3296 3677 -3262 3695
rect -2854 5565 -2820 5583
rect -2854 5549 -2820 5565
rect -2854 5497 -2820 5511
rect -2854 5477 -2820 5497
rect -2854 5429 -2820 5439
rect -2854 5405 -2820 5429
rect -2854 5361 -2820 5367
rect -2854 5333 -2820 5361
rect -2854 5293 -2820 5295
rect -2854 5261 -2820 5293
rect -2854 5191 -2820 5223
rect -2854 5189 -2820 5191
rect -2854 5123 -2820 5151
rect -2854 5117 -2820 5123
rect -2854 5055 -2820 5079
rect -2854 5045 -2820 5055
rect -2854 4987 -2820 5007
rect -2854 4973 -2820 4987
rect -2854 4919 -2820 4935
rect -2854 4901 -2820 4919
rect -2854 4851 -2820 4863
rect -2854 4829 -2820 4851
rect -2854 4783 -2820 4791
rect -2854 4757 -2820 4783
rect -2854 4715 -2820 4719
rect -2854 4685 -2820 4715
rect -2854 4613 -2820 4647
rect -2854 4545 -2820 4575
rect -2854 4541 -2820 4545
rect -2854 4477 -2820 4503
rect -2854 4469 -2820 4477
rect -2854 4409 -2820 4431
rect -2854 4397 -2820 4409
rect -2854 4341 -2820 4359
rect -2854 4325 -2820 4341
rect -2854 4273 -2820 4287
rect -2854 4253 -2820 4273
rect -2854 4205 -2820 4215
rect -2854 4181 -2820 4205
rect -2854 4137 -2820 4143
rect -2854 4109 -2820 4137
rect -2854 4069 -2820 4071
rect -2854 4037 -2820 4069
rect -2854 3967 -2820 3999
rect -2854 3965 -2820 3967
rect -2854 3899 -2820 3927
rect -2854 3893 -2820 3899
rect -2854 3831 -2820 3855
rect -2854 3821 -2820 3831
rect -2854 3763 -2820 3783
rect -2854 3749 -2820 3763
rect -2854 3695 -2820 3711
rect -2854 3677 -2820 3695
rect -2596 5565 -2562 5583
rect -2596 5549 -2562 5565
rect -2596 5497 -2562 5511
rect -2596 5477 -2562 5497
rect -2596 5429 -2562 5439
rect -2596 5405 -2562 5429
rect -2596 5361 -2562 5367
rect -2596 5333 -2562 5361
rect -2596 5293 -2562 5295
rect -2596 5261 -2562 5293
rect -2596 5191 -2562 5223
rect -2596 5189 -2562 5191
rect -2596 5123 -2562 5151
rect -2596 5117 -2562 5123
rect -2596 5055 -2562 5079
rect -2596 5045 -2562 5055
rect -2596 4987 -2562 5007
rect -2596 4973 -2562 4987
rect -2596 4919 -2562 4935
rect -2596 4901 -2562 4919
rect -2596 4851 -2562 4863
rect -2596 4829 -2562 4851
rect -2596 4783 -2562 4791
rect -2596 4757 -2562 4783
rect -2596 4715 -2562 4719
rect -2596 4685 -2562 4715
rect -2596 4613 -2562 4647
rect -2596 4545 -2562 4575
rect -2596 4541 -2562 4545
rect -2596 4477 -2562 4503
rect -2596 4469 -2562 4477
rect -2596 4409 -2562 4431
rect -2596 4397 -2562 4409
rect -2596 4341 -2562 4359
rect -2596 4325 -2562 4341
rect -2596 4273 -2562 4287
rect -2596 4253 -2562 4273
rect -2596 4205 -2562 4215
rect -2596 4181 -2562 4205
rect -2596 4137 -2562 4143
rect -2596 4109 -2562 4137
rect -2596 4069 -2562 4071
rect -2596 4037 -2562 4069
rect -2596 3967 -2562 3999
rect -2596 3965 -2562 3967
rect -2596 3899 -2562 3927
rect -2596 3893 -2562 3899
rect -2596 3831 -2562 3855
rect -2596 3821 -2562 3831
rect -2596 3763 -2562 3783
rect -2596 3749 -2562 3763
rect -2596 3695 -2562 3711
rect -2596 3677 -2562 3695
rect -2154 5565 -2120 5583
rect -2154 5549 -2120 5565
rect -2154 5497 -2120 5511
rect -2154 5477 -2120 5497
rect -2154 5429 -2120 5439
rect -2154 5405 -2120 5429
rect -2154 5361 -2120 5367
rect -2154 5333 -2120 5361
rect -2154 5293 -2120 5295
rect -2154 5261 -2120 5293
rect -2154 5191 -2120 5223
rect -2154 5189 -2120 5191
rect -2154 5123 -2120 5151
rect -2154 5117 -2120 5123
rect -2154 5055 -2120 5079
rect -2154 5045 -2120 5055
rect -2154 4987 -2120 5007
rect -2154 4973 -2120 4987
rect -2154 4919 -2120 4935
rect -2154 4901 -2120 4919
rect -2154 4851 -2120 4863
rect -2154 4829 -2120 4851
rect -2154 4783 -2120 4791
rect -2154 4757 -2120 4783
rect -2154 4715 -2120 4719
rect -2154 4685 -2120 4715
rect -2154 4613 -2120 4647
rect -2154 4545 -2120 4575
rect -2154 4541 -2120 4545
rect -2154 4477 -2120 4503
rect -2154 4469 -2120 4477
rect -2154 4409 -2120 4431
rect -2154 4397 -2120 4409
rect -2154 4341 -2120 4359
rect -2154 4325 -2120 4341
rect -2154 4273 -2120 4287
rect -2154 4253 -2120 4273
rect -2154 4205 -2120 4215
rect -2154 4181 -2120 4205
rect -2154 4137 -2120 4143
rect -2154 4109 -2120 4137
rect -2154 4069 -2120 4071
rect -2154 4037 -2120 4069
rect -2154 3967 -2120 3999
rect -2154 3965 -2120 3967
rect -2154 3899 -2120 3927
rect -2154 3893 -2120 3899
rect -2154 3831 -2120 3855
rect -2154 3821 -2120 3831
rect -2154 3763 -2120 3783
rect -2154 3749 -2120 3763
rect -2154 3695 -2120 3711
rect -2154 3677 -2120 3695
rect -1896 5565 -1862 5583
rect -1896 5549 -1862 5565
rect -1896 5497 -1862 5511
rect -1896 5477 -1862 5497
rect -1896 5429 -1862 5439
rect -1896 5405 -1862 5429
rect -1896 5361 -1862 5367
rect -1896 5333 -1862 5361
rect -1896 5293 -1862 5295
rect -1896 5261 -1862 5293
rect -1896 5191 -1862 5223
rect -1896 5189 -1862 5191
rect -1896 5123 -1862 5151
rect -1896 5117 -1862 5123
rect -1896 5055 -1862 5079
rect -1896 5045 -1862 5055
rect -1896 4987 -1862 5007
rect -1896 4973 -1862 4987
rect -1896 4919 -1862 4935
rect -1896 4901 -1862 4919
rect -1896 4851 -1862 4863
rect -1896 4829 -1862 4851
rect -1896 4783 -1862 4791
rect -1896 4757 -1862 4783
rect -1896 4715 -1862 4719
rect -1896 4685 -1862 4715
rect -1896 4613 -1862 4647
rect -1896 4545 -1862 4575
rect -1896 4541 -1862 4545
rect -1896 4477 -1862 4503
rect -1896 4469 -1862 4477
rect -1896 4409 -1862 4431
rect -1896 4397 -1862 4409
rect -1896 4341 -1862 4359
rect -1896 4325 -1862 4341
rect -1896 4273 -1862 4287
rect -1896 4253 -1862 4273
rect -1896 4205 -1862 4215
rect -1896 4181 -1862 4205
rect -1896 4137 -1862 4143
rect -1896 4109 -1862 4137
rect -1896 4069 -1862 4071
rect -1896 4037 -1862 4069
rect -1896 3967 -1862 3999
rect -1896 3965 -1862 3967
rect -1896 3899 -1862 3927
rect -1896 3893 -1862 3899
rect -1896 3831 -1862 3855
rect -1896 3821 -1862 3831
rect -1896 3763 -1862 3783
rect -1896 3749 -1862 3763
rect -1896 3695 -1862 3711
rect -1896 3677 -1862 3695
rect -1454 5565 -1420 5583
rect -1454 5549 -1420 5565
rect -1454 5497 -1420 5511
rect -1454 5477 -1420 5497
rect -1454 5429 -1420 5439
rect -1454 5405 -1420 5429
rect -1454 5361 -1420 5367
rect -1454 5333 -1420 5361
rect -1454 5293 -1420 5295
rect -1454 5261 -1420 5293
rect -1454 5191 -1420 5223
rect -1454 5189 -1420 5191
rect -1454 5123 -1420 5151
rect -1454 5117 -1420 5123
rect -1454 5055 -1420 5079
rect -1454 5045 -1420 5055
rect -1454 4987 -1420 5007
rect -1454 4973 -1420 4987
rect -1454 4919 -1420 4935
rect -1454 4901 -1420 4919
rect -1454 4851 -1420 4863
rect -1454 4829 -1420 4851
rect -1454 4783 -1420 4791
rect -1454 4757 -1420 4783
rect -1454 4715 -1420 4719
rect -1454 4685 -1420 4715
rect -1454 4613 -1420 4647
rect -1454 4545 -1420 4575
rect -1454 4541 -1420 4545
rect -1454 4477 -1420 4503
rect -1454 4469 -1420 4477
rect -1454 4409 -1420 4431
rect -1454 4397 -1420 4409
rect -1454 4341 -1420 4359
rect -1454 4325 -1420 4341
rect -1454 4273 -1420 4287
rect -1454 4253 -1420 4273
rect -1454 4205 -1420 4215
rect -1454 4181 -1420 4205
rect -1454 4137 -1420 4143
rect -1454 4109 -1420 4137
rect -1454 4069 -1420 4071
rect -1454 4037 -1420 4069
rect -1454 3967 -1420 3999
rect -1454 3965 -1420 3967
rect -1454 3899 -1420 3927
rect -1454 3893 -1420 3899
rect -1454 3831 -1420 3855
rect -1454 3821 -1420 3831
rect -1454 3763 -1420 3783
rect -1454 3749 -1420 3763
rect -1454 3695 -1420 3711
rect -1454 3677 -1420 3695
rect -1196 5565 -1162 5583
rect -1196 5549 -1162 5565
rect -1196 5497 -1162 5511
rect -1196 5477 -1162 5497
rect -1196 5429 -1162 5439
rect -1196 5405 -1162 5429
rect -1196 5361 -1162 5367
rect -1196 5333 -1162 5361
rect -1196 5293 -1162 5295
rect -1196 5261 -1162 5293
rect -1196 5191 -1162 5223
rect -1196 5189 -1162 5191
rect -1196 5123 -1162 5151
rect -1196 5117 -1162 5123
rect -1196 5055 -1162 5079
rect -1196 5045 -1162 5055
rect -1196 4987 -1162 5007
rect -1196 4973 -1162 4987
rect -1196 4919 -1162 4935
rect -1196 4901 -1162 4919
rect -1196 4851 -1162 4863
rect -1196 4829 -1162 4851
rect -1196 4783 -1162 4791
rect -1196 4757 -1162 4783
rect -1196 4715 -1162 4719
rect -1196 4685 -1162 4715
rect -1196 4613 -1162 4647
rect -1196 4545 -1162 4575
rect -1196 4541 -1162 4545
rect -1196 4477 -1162 4503
rect -1196 4469 -1162 4477
rect -1196 4409 -1162 4431
rect -1196 4397 -1162 4409
rect -1196 4341 -1162 4359
rect -1196 4325 -1162 4341
rect -1196 4273 -1162 4287
rect -1196 4253 -1162 4273
rect -1196 4205 -1162 4215
rect -1196 4181 -1162 4205
rect -1196 4137 -1162 4143
rect -1196 4109 -1162 4137
rect -1196 4069 -1162 4071
rect -1196 4037 -1162 4069
rect -1196 3967 -1162 3999
rect -1196 3965 -1162 3967
rect -1196 3899 -1162 3927
rect -1196 3893 -1162 3899
rect -1196 3831 -1162 3855
rect -1196 3821 -1162 3831
rect -1196 3763 -1162 3783
rect -1196 3749 -1162 3763
rect -1196 3695 -1162 3711
rect -1196 3677 -1162 3695
rect -754 5565 -720 5583
rect -754 5549 -720 5565
rect -754 5497 -720 5511
rect -754 5477 -720 5497
rect -754 5429 -720 5439
rect -754 5405 -720 5429
rect -754 5361 -720 5367
rect -754 5333 -720 5361
rect -754 5293 -720 5295
rect -754 5261 -720 5293
rect -754 5191 -720 5223
rect -754 5189 -720 5191
rect -754 5123 -720 5151
rect -754 5117 -720 5123
rect -754 5055 -720 5079
rect -754 5045 -720 5055
rect -754 4987 -720 5007
rect -754 4973 -720 4987
rect -754 4919 -720 4935
rect -754 4901 -720 4919
rect -754 4851 -720 4863
rect -754 4829 -720 4851
rect -754 4783 -720 4791
rect -754 4757 -720 4783
rect -754 4715 -720 4719
rect -754 4685 -720 4715
rect -754 4613 -720 4647
rect -754 4545 -720 4575
rect -754 4541 -720 4545
rect -754 4477 -720 4503
rect -754 4469 -720 4477
rect -754 4409 -720 4431
rect -754 4397 -720 4409
rect -754 4341 -720 4359
rect -754 4325 -720 4341
rect -754 4273 -720 4287
rect -754 4253 -720 4273
rect -754 4205 -720 4215
rect -754 4181 -720 4205
rect -754 4137 -720 4143
rect -754 4109 -720 4137
rect -754 4069 -720 4071
rect -754 4037 -720 4069
rect -754 3967 -720 3999
rect -754 3965 -720 3967
rect -754 3899 -720 3927
rect -754 3893 -720 3899
rect -754 3831 -720 3855
rect -754 3821 -720 3831
rect -754 3763 -720 3783
rect -754 3749 -720 3763
rect -754 3695 -720 3711
rect -754 3677 -720 3695
rect -496 5565 -462 5583
rect -496 5549 -462 5565
rect -496 5497 -462 5511
rect -496 5477 -462 5497
rect -496 5429 -462 5439
rect -496 5405 -462 5429
rect -496 5361 -462 5367
rect -496 5333 -462 5361
rect -496 5293 -462 5295
rect -496 5261 -462 5293
rect -496 5191 -462 5223
rect -496 5189 -462 5191
rect -496 5123 -462 5151
rect -496 5117 -462 5123
rect -496 5055 -462 5079
rect -496 5045 -462 5055
rect -496 4987 -462 5007
rect -496 4973 -462 4987
rect -496 4919 -462 4935
rect -496 4901 -462 4919
rect -496 4851 -462 4863
rect -496 4829 -462 4851
rect -496 4783 -462 4791
rect -496 4757 -462 4783
rect -496 4715 -462 4719
rect -496 4685 -462 4715
rect -496 4613 -462 4647
rect -496 4545 -462 4575
rect -496 4541 -462 4545
rect -496 4477 -462 4503
rect -496 4469 -462 4477
rect -496 4409 -462 4431
rect -496 4397 -462 4409
rect -496 4341 -462 4359
rect -496 4325 -462 4341
rect -496 4273 -462 4287
rect -496 4253 -462 4273
rect -496 4205 -462 4215
rect -496 4181 -462 4205
rect -496 4137 -462 4143
rect -496 4109 -462 4137
rect -496 4069 -462 4071
rect -496 4037 -462 4069
rect -496 3967 -462 3999
rect -496 3965 -462 3967
rect -496 3899 -462 3927
rect -496 3893 -462 3899
rect -496 3831 -462 3855
rect -496 3821 -462 3831
rect -496 3763 -462 3783
rect -496 3749 -462 3763
rect -496 3695 -462 3711
rect -496 3677 -462 3695
rect -54 5565 -20 5583
rect -54 5549 -20 5565
rect -54 5497 -20 5511
rect -54 5477 -20 5497
rect -54 5429 -20 5439
rect -54 5405 -20 5429
rect -54 5361 -20 5367
rect -54 5333 -20 5361
rect -54 5293 -20 5295
rect -54 5261 -20 5293
rect -54 5191 -20 5223
rect -54 5189 -20 5191
rect -54 5123 -20 5151
rect -54 5117 -20 5123
rect -54 5055 -20 5079
rect -54 5045 -20 5055
rect -54 4987 -20 5007
rect -54 4973 -20 4987
rect -54 4919 -20 4935
rect -54 4901 -20 4919
rect -54 4851 -20 4863
rect -54 4829 -20 4851
rect -54 4783 -20 4791
rect -54 4757 -20 4783
rect -54 4715 -20 4719
rect -54 4685 -20 4715
rect -54 4613 -20 4647
rect -54 4545 -20 4575
rect -54 4541 -20 4545
rect -54 4477 -20 4503
rect -54 4469 -20 4477
rect -54 4409 -20 4431
rect -54 4397 -20 4409
rect -54 4341 -20 4359
rect -54 4325 -20 4341
rect -54 4273 -20 4287
rect -54 4253 -20 4273
rect -54 4205 -20 4215
rect -54 4181 -20 4205
rect -54 4137 -20 4143
rect -54 4109 -20 4137
rect -54 4069 -20 4071
rect -54 4037 -20 4069
rect -54 3967 -20 3999
rect -54 3965 -20 3967
rect -54 3899 -20 3927
rect -54 3893 -20 3899
rect -54 3831 -20 3855
rect -54 3821 -20 3831
rect -54 3763 -20 3783
rect -54 3749 -20 3763
rect -54 3695 -20 3711
rect -54 3677 -20 3695
rect 204 5565 238 5583
rect 204 5549 238 5565
rect 204 5497 238 5511
rect 204 5477 238 5497
rect 204 5429 238 5439
rect 204 5405 238 5429
rect 204 5361 238 5367
rect 204 5333 238 5361
rect 204 5293 238 5295
rect 204 5261 238 5293
rect 204 5191 238 5223
rect 204 5189 238 5191
rect 204 5123 238 5151
rect 204 5117 238 5123
rect 204 5055 238 5079
rect 204 5045 238 5055
rect 204 4987 238 5007
rect 204 4973 238 4987
rect 204 4919 238 4935
rect 204 4901 238 4919
rect 204 4851 238 4863
rect 204 4829 238 4851
rect 204 4783 238 4791
rect 204 4757 238 4783
rect 204 4715 238 4719
rect 204 4685 238 4715
rect 204 4613 238 4647
rect 204 4545 238 4575
rect 204 4541 238 4545
rect 204 4477 238 4503
rect 204 4469 238 4477
rect 204 4409 238 4431
rect 204 4397 238 4409
rect 204 4341 238 4359
rect 204 4325 238 4341
rect 204 4273 238 4287
rect 204 4253 238 4273
rect 204 4205 238 4215
rect 204 4181 238 4205
rect 204 4137 238 4143
rect 204 4109 238 4137
rect 204 4069 238 4071
rect 204 4037 238 4069
rect 204 3967 238 3999
rect 204 3965 238 3967
rect 204 3899 238 3927
rect 204 3893 238 3899
rect 204 3831 238 3855
rect 204 3821 238 3831
rect 204 3763 238 3783
rect 204 3749 238 3763
rect 204 3695 238 3711
rect 204 3677 238 3695
rect 646 5565 680 5583
rect 646 5549 680 5565
rect 646 5497 680 5511
rect 646 5477 680 5497
rect 646 5429 680 5439
rect 646 5405 680 5429
rect 646 5361 680 5367
rect 646 5333 680 5361
rect 646 5293 680 5295
rect 646 5261 680 5293
rect 646 5191 680 5223
rect 646 5189 680 5191
rect 646 5123 680 5151
rect 646 5117 680 5123
rect 646 5055 680 5079
rect 646 5045 680 5055
rect 646 4987 680 5007
rect 646 4973 680 4987
rect 646 4919 680 4935
rect 646 4901 680 4919
rect 646 4851 680 4863
rect 646 4829 680 4851
rect 646 4783 680 4791
rect 646 4757 680 4783
rect 646 4715 680 4719
rect 646 4685 680 4715
rect 646 4613 680 4647
rect 646 4545 680 4575
rect 646 4541 680 4545
rect 646 4477 680 4503
rect 646 4469 680 4477
rect 646 4409 680 4431
rect 646 4397 680 4409
rect 646 4341 680 4359
rect 646 4325 680 4341
rect 646 4273 680 4287
rect 646 4253 680 4273
rect 646 4205 680 4215
rect 646 4181 680 4205
rect 646 4137 680 4143
rect 646 4109 680 4137
rect 646 4069 680 4071
rect 646 4037 680 4069
rect 646 3967 680 3999
rect 646 3965 680 3967
rect 646 3899 680 3927
rect 646 3893 680 3899
rect 646 3831 680 3855
rect 646 3821 680 3831
rect 646 3763 680 3783
rect 646 3749 680 3763
rect 646 3695 680 3711
rect 646 3677 680 3695
rect 904 5565 938 5583
rect 904 5549 938 5565
rect 904 5497 938 5511
rect 904 5477 938 5497
rect 904 5429 938 5439
rect 904 5405 938 5429
rect 904 5361 938 5367
rect 904 5333 938 5361
rect 904 5293 938 5295
rect 904 5261 938 5293
rect 904 5191 938 5223
rect 904 5189 938 5191
rect 904 5123 938 5151
rect 904 5117 938 5123
rect 904 5055 938 5079
rect 904 5045 938 5055
rect 904 4987 938 5007
rect 904 4973 938 4987
rect 904 4919 938 4935
rect 904 4901 938 4919
rect 904 4851 938 4863
rect 904 4829 938 4851
rect 904 4783 938 4791
rect 904 4757 938 4783
rect 904 4715 938 4719
rect 904 4685 938 4715
rect 904 4613 938 4647
rect 904 4545 938 4575
rect 904 4541 938 4545
rect 904 4477 938 4503
rect 904 4469 938 4477
rect 904 4409 938 4431
rect 904 4397 938 4409
rect 904 4341 938 4359
rect 904 4325 938 4341
rect 904 4273 938 4287
rect 904 4253 938 4273
rect 904 4205 938 4215
rect 904 4181 938 4205
rect 904 4137 938 4143
rect 904 4109 938 4137
rect 904 4069 938 4071
rect 904 4037 938 4069
rect 904 3967 938 3999
rect 904 3965 938 3967
rect 904 3899 938 3927
rect 904 3893 938 3899
rect 904 3831 938 3855
rect 904 3821 938 3831
rect 904 3763 938 3783
rect 904 3749 938 3763
rect 904 3695 938 3711
rect 904 3677 938 3695
rect 1346 5565 1380 5583
rect 1346 5549 1380 5565
rect 1346 5497 1380 5511
rect 1346 5477 1380 5497
rect 1346 5429 1380 5439
rect 1346 5405 1380 5429
rect 1346 5361 1380 5367
rect 1346 5333 1380 5361
rect 1346 5293 1380 5295
rect 1346 5261 1380 5293
rect 1346 5191 1380 5223
rect 1346 5189 1380 5191
rect 1346 5123 1380 5151
rect 1346 5117 1380 5123
rect 1346 5055 1380 5079
rect 1346 5045 1380 5055
rect 1346 4987 1380 5007
rect 1346 4973 1380 4987
rect 1346 4919 1380 4935
rect 1346 4901 1380 4919
rect 1346 4851 1380 4863
rect 1346 4829 1380 4851
rect 1346 4783 1380 4791
rect 1346 4757 1380 4783
rect 1346 4715 1380 4719
rect 1346 4685 1380 4715
rect 1346 4613 1380 4647
rect 1346 4545 1380 4575
rect 1346 4541 1380 4545
rect 1346 4477 1380 4503
rect 1346 4469 1380 4477
rect 1346 4409 1380 4431
rect 1346 4397 1380 4409
rect 1346 4341 1380 4359
rect 1346 4325 1380 4341
rect 1346 4273 1380 4287
rect 1346 4253 1380 4273
rect 1346 4205 1380 4215
rect 1346 4181 1380 4205
rect 1346 4137 1380 4143
rect 1346 4109 1380 4137
rect 1346 4069 1380 4071
rect 1346 4037 1380 4069
rect 1346 3967 1380 3999
rect 1346 3965 1380 3967
rect 1346 3899 1380 3927
rect 1346 3893 1380 3899
rect 1346 3831 1380 3855
rect 1346 3821 1380 3831
rect 1346 3763 1380 3783
rect 1346 3749 1380 3763
rect 1346 3695 1380 3711
rect 1346 3677 1380 3695
rect 1604 5565 1638 5583
rect 1604 5549 1638 5565
rect 1604 5497 1638 5511
rect 1604 5477 1638 5497
rect 1604 5429 1638 5439
rect 1604 5405 1638 5429
rect 1604 5361 1638 5367
rect 1604 5333 1638 5361
rect 1604 5293 1638 5295
rect 1604 5261 1638 5293
rect 1604 5191 1638 5223
rect 1604 5189 1638 5191
rect 1604 5123 1638 5151
rect 1604 5117 1638 5123
rect 1604 5055 1638 5079
rect 1604 5045 1638 5055
rect 1604 4987 1638 5007
rect 1604 4973 1638 4987
rect 1604 4919 1638 4935
rect 1604 4901 1638 4919
rect 1604 4851 1638 4863
rect 1604 4829 1638 4851
rect 1604 4783 1638 4791
rect 1604 4757 1638 4783
rect 1604 4715 1638 4719
rect 1604 4685 1638 4715
rect 1604 4613 1638 4647
rect 1604 4545 1638 4575
rect 1604 4541 1638 4545
rect 1604 4477 1638 4503
rect 1604 4469 1638 4477
rect 1604 4409 1638 4431
rect 1604 4397 1638 4409
rect 1604 4341 1638 4359
rect 1604 4325 1638 4341
rect 1604 4273 1638 4287
rect 1604 4253 1638 4273
rect 1604 4205 1638 4215
rect 1604 4181 1638 4205
rect 1604 4137 1638 4143
rect 1604 4109 1638 4137
rect 1604 4069 1638 4071
rect 1604 4037 1638 4069
rect 1604 3967 1638 3999
rect 1604 3965 1638 3967
rect 1604 3899 1638 3927
rect 1604 3893 1638 3899
rect 1604 3831 1638 3855
rect 1604 3821 1638 3831
rect 1604 3763 1638 3783
rect 1604 3749 1638 3763
rect 1604 3695 1638 3711
rect 1604 3677 1638 3695
rect 2046 5565 2080 5583
rect 2046 5549 2080 5565
rect 2046 5497 2080 5511
rect 2046 5477 2080 5497
rect 2046 5429 2080 5439
rect 2046 5405 2080 5429
rect 2046 5361 2080 5367
rect 2046 5333 2080 5361
rect 2046 5293 2080 5295
rect 2046 5261 2080 5293
rect 2046 5191 2080 5223
rect 2046 5189 2080 5191
rect 2046 5123 2080 5151
rect 2046 5117 2080 5123
rect 2046 5055 2080 5079
rect 2046 5045 2080 5055
rect 2046 4987 2080 5007
rect 2046 4973 2080 4987
rect 2046 4919 2080 4935
rect 2046 4901 2080 4919
rect 2046 4851 2080 4863
rect 2046 4829 2080 4851
rect 2046 4783 2080 4791
rect 2046 4757 2080 4783
rect 2046 4715 2080 4719
rect 2046 4685 2080 4715
rect 2046 4613 2080 4647
rect 2046 4545 2080 4575
rect 2046 4541 2080 4545
rect 2046 4477 2080 4503
rect 2046 4469 2080 4477
rect 2046 4409 2080 4431
rect 2046 4397 2080 4409
rect 2046 4341 2080 4359
rect 2046 4325 2080 4341
rect 2046 4273 2080 4287
rect 2046 4253 2080 4273
rect 2046 4205 2080 4215
rect 2046 4181 2080 4205
rect 2046 4137 2080 4143
rect 2046 4109 2080 4137
rect 2046 4069 2080 4071
rect 2046 4037 2080 4069
rect 2046 3967 2080 3999
rect 2046 3965 2080 3967
rect 2046 3899 2080 3927
rect 2046 3893 2080 3899
rect 2046 3831 2080 3855
rect 2046 3821 2080 3831
rect 2046 3763 2080 3783
rect 2046 3749 2080 3763
rect 2046 3695 2080 3711
rect 2046 3677 2080 3695
rect 2304 5565 2338 5583
rect 2304 5549 2338 5565
rect 2304 5497 2338 5511
rect 2304 5477 2338 5497
rect 2304 5429 2338 5439
rect 2304 5405 2338 5429
rect 2304 5361 2338 5367
rect 2304 5333 2338 5361
rect 2304 5293 2338 5295
rect 2304 5261 2338 5293
rect 2304 5191 2338 5223
rect 2304 5189 2338 5191
rect 2304 5123 2338 5151
rect 2304 5117 2338 5123
rect 2304 5055 2338 5079
rect 2304 5045 2338 5055
rect 2304 4987 2338 5007
rect 2304 4973 2338 4987
rect 2304 4919 2338 4935
rect 2304 4901 2338 4919
rect 2304 4851 2338 4863
rect 2304 4829 2338 4851
rect 2304 4783 2338 4791
rect 2304 4757 2338 4783
rect 2304 4715 2338 4719
rect 2304 4685 2338 4715
rect 2304 4613 2338 4647
rect 2304 4545 2338 4575
rect 2304 4541 2338 4545
rect 2304 4477 2338 4503
rect 2304 4469 2338 4477
rect 2304 4409 2338 4431
rect 2304 4397 2338 4409
rect 2304 4341 2338 4359
rect 2304 4325 2338 4341
rect 2304 4273 2338 4287
rect 2304 4253 2338 4273
rect 2304 4205 2338 4215
rect 2304 4181 2338 4205
rect 2304 4137 2338 4143
rect 2304 4109 2338 4137
rect 2304 4069 2338 4071
rect 2304 4037 2338 4069
rect 2304 3967 2338 3999
rect 2304 3965 2338 3967
rect 2304 3899 2338 3927
rect 2304 3893 2338 3899
rect 2304 3831 2338 3855
rect 2304 3821 2338 3831
rect 2304 3763 2338 3783
rect 2304 3749 2338 3763
rect 2304 3695 2338 3711
rect 2304 3677 2338 3695
rect 3746 5565 3780 5583
rect 3746 5549 3780 5565
rect 3746 5497 3780 5511
rect 3746 5477 3780 5497
rect 3746 5429 3780 5439
rect 3746 5405 3780 5429
rect 3746 5361 3780 5367
rect 3746 5333 3780 5361
rect 3746 5293 3780 5295
rect 3746 5261 3780 5293
rect 3746 5191 3780 5223
rect 3746 5189 3780 5191
rect 3746 5123 3780 5151
rect 3746 5117 3780 5123
rect 3746 5055 3780 5079
rect 3746 5045 3780 5055
rect 3746 4987 3780 5007
rect 3746 4973 3780 4987
rect 3746 4919 3780 4935
rect 3746 4901 3780 4919
rect 3746 4851 3780 4863
rect 3746 4829 3780 4851
rect 3746 4783 3780 4791
rect 3746 4757 3780 4783
rect 3746 4715 3780 4719
rect 3746 4685 3780 4715
rect 3746 4613 3780 4647
rect 3746 4545 3780 4575
rect 3746 4541 3780 4545
rect 3746 4477 3780 4503
rect 3746 4469 3780 4477
rect 3746 4409 3780 4431
rect 3746 4397 3780 4409
rect 3746 4341 3780 4359
rect 3746 4325 3780 4341
rect 3746 4273 3780 4287
rect 3746 4253 3780 4273
rect 3746 4205 3780 4215
rect 3746 4181 3780 4205
rect 3746 4137 3780 4143
rect 3746 4109 3780 4137
rect 3746 4069 3780 4071
rect 3746 4037 3780 4069
rect 3746 3967 3780 3999
rect 3746 3965 3780 3967
rect 3746 3899 3780 3927
rect 3746 3893 3780 3899
rect 3746 3831 3780 3855
rect 3746 3821 3780 3831
rect 3746 3763 3780 3783
rect 3746 3749 3780 3763
rect 3746 3695 3780 3711
rect 3746 3677 3780 3695
rect 4004 5565 4038 5583
rect 4004 5549 4038 5565
rect 4004 5497 4038 5511
rect 4004 5477 4038 5497
rect 4004 5429 4038 5439
rect 4004 5405 4038 5429
rect 4004 5361 4038 5367
rect 4004 5333 4038 5361
rect 4004 5293 4038 5295
rect 4004 5261 4038 5293
rect 4004 5191 4038 5223
rect 4004 5189 4038 5191
rect 4004 5123 4038 5151
rect 4004 5117 4038 5123
rect 4004 5055 4038 5079
rect 4004 5045 4038 5055
rect 4004 4987 4038 5007
rect 4004 4973 4038 4987
rect 4004 4919 4038 4935
rect 4004 4901 4038 4919
rect 4004 4851 4038 4863
rect 4004 4829 4038 4851
rect 4004 4783 4038 4791
rect 4004 4757 4038 4783
rect 4004 4715 4038 4719
rect 4004 4685 4038 4715
rect 4004 4613 4038 4647
rect 4004 4545 4038 4575
rect 4004 4541 4038 4545
rect 4004 4477 4038 4503
rect 4004 4469 4038 4477
rect 4004 4409 4038 4431
rect 4004 4397 4038 4409
rect 4004 4341 4038 4359
rect 4004 4325 4038 4341
rect 4004 4273 4038 4287
rect 4004 4253 4038 4273
rect 4004 4205 4038 4215
rect 4004 4181 4038 4205
rect 4004 4137 4038 4143
rect 4004 4109 4038 4137
rect 4004 4069 4038 4071
rect 4004 4037 4038 4069
rect 4004 3967 4038 3999
rect 4004 3965 4038 3967
rect 4004 3899 4038 3927
rect 4004 3893 4038 3899
rect 4004 3831 4038 3855
rect 4004 3821 4038 3831
rect 4004 3763 4038 3783
rect 4004 3749 4038 3763
rect 4004 3695 4038 3711
rect 4004 3677 4038 3695
rect 4446 5565 4480 5583
rect 4446 5549 4480 5565
rect 4446 5497 4480 5511
rect 4446 5477 4480 5497
rect 4446 5429 4480 5439
rect 4446 5405 4480 5429
rect 4446 5361 4480 5367
rect 4446 5333 4480 5361
rect 4446 5293 4480 5295
rect 4446 5261 4480 5293
rect 4446 5191 4480 5223
rect 4446 5189 4480 5191
rect 4446 5123 4480 5151
rect 4446 5117 4480 5123
rect 4446 5055 4480 5079
rect 4446 5045 4480 5055
rect 4446 4987 4480 5007
rect 4446 4973 4480 4987
rect 4446 4919 4480 4935
rect 4446 4901 4480 4919
rect 4446 4851 4480 4863
rect 4446 4829 4480 4851
rect 4446 4783 4480 4791
rect 4446 4757 4480 4783
rect 4446 4715 4480 4719
rect 4446 4685 4480 4715
rect 4446 4613 4480 4647
rect 4446 4545 4480 4575
rect 4446 4541 4480 4545
rect 4446 4477 4480 4503
rect 4446 4469 4480 4477
rect 4446 4409 4480 4431
rect 4446 4397 4480 4409
rect 4446 4341 4480 4359
rect 4446 4325 4480 4341
rect 4446 4273 4480 4287
rect 4446 4253 4480 4273
rect 4446 4205 4480 4215
rect 4446 4181 4480 4205
rect 4446 4137 4480 4143
rect 4446 4109 4480 4137
rect 4446 4069 4480 4071
rect 4446 4037 4480 4069
rect 4446 3967 4480 3999
rect 4446 3965 4480 3967
rect 4446 3899 4480 3927
rect 4446 3893 4480 3899
rect 4446 3831 4480 3855
rect 4446 3821 4480 3831
rect 4446 3763 4480 3783
rect 4446 3749 4480 3763
rect 4446 3695 4480 3711
rect 4446 3677 4480 3695
rect 4704 5565 4738 5583
rect 4704 5549 4738 5565
rect 4704 5497 4738 5511
rect 4704 5477 4738 5497
rect 4704 5429 4738 5439
rect 4704 5405 4738 5429
rect 4704 5361 4738 5367
rect 4704 5333 4738 5361
rect 4704 5293 4738 5295
rect 4704 5261 4738 5293
rect 4704 5191 4738 5223
rect 4704 5189 4738 5191
rect 4704 5123 4738 5151
rect 4704 5117 4738 5123
rect 4704 5055 4738 5079
rect 4704 5045 4738 5055
rect 4704 4987 4738 5007
rect 4704 4973 4738 4987
rect 4704 4919 4738 4935
rect 4704 4901 4738 4919
rect 4704 4851 4738 4863
rect 4704 4829 4738 4851
rect 4704 4783 4738 4791
rect 4704 4757 4738 4783
rect 4704 4715 4738 4719
rect 4704 4685 4738 4715
rect 4704 4613 4738 4647
rect 4704 4545 4738 4575
rect 4704 4541 4738 4545
rect 4704 4477 4738 4503
rect 4704 4469 4738 4477
rect 4704 4409 4738 4431
rect 4704 4397 4738 4409
rect 4704 4341 4738 4359
rect 4704 4325 4738 4341
rect 4704 4273 4738 4287
rect 4704 4253 4738 4273
rect 4704 4205 4738 4215
rect 4704 4181 4738 4205
rect 4704 4137 4738 4143
rect 4704 4109 4738 4137
rect 4704 4069 4738 4071
rect 4704 4037 4738 4069
rect 4704 3967 4738 3999
rect 4704 3965 4738 3967
rect 4704 3899 4738 3927
rect 4704 3893 4738 3899
rect 4704 3831 4738 3855
rect 4704 3821 4738 3831
rect 4704 3763 4738 3783
rect 4704 3749 4738 3763
rect 4704 3695 4738 3711
rect 4704 3677 4738 3695
rect 5146 5565 5180 5583
rect 5146 5549 5180 5565
rect 5146 5497 5180 5511
rect 5146 5477 5180 5497
rect 5146 5429 5180 5439
rect 5146 5405 5180 5429
rect 5146 5361 5180 5367
rect 5146 5333 5180 5361
rect 5146 5293 5180 5295
rect 5146 5261 5180 5293
rect 5146 5191 5180 5223
rect 5146 5189 5180 5191
rect 5146 5123 5180 5151
rect 5146 5117 5180 5123
rect 5146 5055 5180 5079
rect 5146 5045 5180 5055
rect 5146 4987 5180 5007
rect 5146 4973 5180 4987
rect 5146 4919 5180 4935
rect 5146 4901 5180 4919
rect 5146 4851 5180 4863
rect 5146 4829 5180 4851
rect 5146 4783 5180 4791
rect 5146 4757 5180 4783
rect 5146 4715 5180 4719
rect 5146 4685 5180 4715
rect 5146 4613 5180 4647
rect 5146 4545 5180 4575
rect 5146 4541 5180 4545
rect 5146 4477 5180 4503
rect 5146 4469 5180 4477
rect 5146 4409 5180 4431
rect 5146 4397 5180 4409
rect 5146 4341 5180 4359
rect 5146 4325 5180 4341
rect 5146 4273 5180 4287
rect 5146 4253 5180 4273
rect 5146 4205 5180 4215
rect 5146 4181 5180 4205
rect 5146 4137 5180 4143
rect 5146 4109 5180 4137
rect 5146 4069 5180 4071
rect 5146 4037 5180 4069
rect 5146 3967 5180 3999
rect 5146 3965 5180 3967
rect 5146 3899 5180 3927
rect 5146 3893 5180 3899
rect 5146 3831 5180 3855
rect 5146 3821 5180 3831
rect 5146 3763 5180 3783
rect 5146 3749 5180 3763
rect 5146 3695 5180 3711
rect 5146 3677 5180 3695
rect 5404 5565 5438 5583
rect 5404 5549 5438 5565
rect 5404 5497 5438 5511
rect 5404 5477 5438 5497
rect 5404 5429 5438 5439
rect 5404 5405 5438 5429
rect 5404 5361 5438 5367
rect 5404 5333 5438 5361
rect 5404 5293 5438 5295
rect 5404 5261 5438 5293
rect 5404 5191 5438 5223
rect 5404 5189 5438 5191
rect 5404 5123 5438 5151
rect 5404 5117 5438 5123
rect 5404 5055 5438 5079
rect 5404 5045 5438 5055
rect 5404 4987 5438 5007
rect 5404 4973 5438 4987
rect 5404 4919 5438 4935
rect 5404 4901 5438 4919
rect 5404 4851 5438 4863
rect 5404 4829 5438 4851
rect 5404 4783 5438 4791
rect 5404 4757 5438 4783
rect 5404 4715 5438 4719
rect 5404 4685 5438 4715
rect 5404 4613 5438 4647
rect 5404 4545 5438 4575
rect 5404 4541 5438 4545
rect 5404 4477 5438 4503
rect 5404 4469 5438 4477
rect 5404 4409 5438 4431
rect 5404 4397 5438 4409
rect 5404 4341 5438 4359
rect 5404 4325 5438 4341
rect 5404 4273 5438 4287
rect 5404 4253 5438 4273
rect 5404 4205 5438 4215
rect 5404 4181 5438 4205
rect 5404 4137 5438 4143
rect 5404 4109 5438 4137
rect 5404 4069 5438 4071
rect 5404 4037 5438 4069
rect 5404 3967 5438 3999
rect 5404 3965 5438 3967
rect 5404 3899 5438 3927
rect 5404 3893 5438 3899
rect 5404 3831 5438 3855
rect 5404 3821 5438 3831
rect 5404 3763 5438 3783
rect 5404 3749 5438 3763
rect 5404 3695 5438 3711
rect 5404 3677 5438 3695
rect 5846 5565 5880 5583
rect 5846 5549 5880 5565
rect 5846 5497 5880 5511
rect 5846 5477 5880 5497
rect 5846 5429 5880 5439
rect 5846 5405 5880 5429
rect 5846 5361 5880 5367
rect 5846 5333 5880 5361
rect 5846 5293 5880 5295
rect 5846 5261 5880 5293
rect 5846 5191 5880 5223
rect 5846 5189 5880 5191
rect 5846 5123 5880 5151
rect 5846 5117 5880 5123
rect 5846 5055 5880 5079
rect 5846 5045 5880 5055
rect 5846 4987 5880 5007
rect 5846 4973 5880 4987
rect 5846 4919 5880 4935
rect 5846 4901 5880 4919
rect 5846 4851 5880 4863
rect 5846 4829 5880 4851
rect 5846 4783 5880 4791
rect 5846 4757 5880 4783
rect 5846 4715 5880 4719
rect 5846 4685 5880 4715
rect 5846 4613 5880 4647
rect 5846 4545 5880 4575
rect 5846 4541 5880 4545
rect 5846 4477 5880 4503
rect 5846 4469 5880 4477
rect 5846 4409 5880 4431
rect 5846 4397 5880 4409
rect 5846 4341 5880 4359
rect 5846 4325 5880 4341
rect 5846 4273 5880 4287
rect 5846 4253 5880 4273
rect 5846 4205 5880 4215
rect 5846 4181 5880 4205
rect 5846 4137 5880 4143
rect 5846 4109 5880 4137
rect 5846 4069 5880 4071
rect 5846 4037 5880 4069
rect 5846 3967 5880 3999
rect 5846 3965 5880 3967
rect 5846 3899 5880 3927
rect 5846 3893 5880 3899
rect 5846 3831 5880 3855
rect 5846 3821 5880 3831
rect 5846 3763 5880 3783
rect 5846 3749 5880 3763
rect 5846 3695 5880 3711
rect 5846 3677 5880 3695
rect 6104 5565 6138 5583
rect 6104 5549 6138 5565
rect 6104 5497 6138 5511
rect 6104 5477 6138 5497
rect 6104 5429 6138 5439
rect 6104 5405 6138 5429
rect 6104 5361 6138 5367
rect 6104 5333 6138 5361
rect 6104 5293 6138 5295
rect 6104 5261 6138 5293
rect 6104 5191 6138 5223
rect 6104 5189 6138 5191
rect 6104 5123 6138 5151
rect 6104 5117 6138 5123
rect 6104 5055 6138 5079
rect 6104 5045 6138 5055
rect 6104 4987 6138 5007
rect 6104 4973 6138 4987
rect 6104 4919 6138 4935
rect 6104 4901 6138 4919
rect 6104 4851 6138 4863
rect 6104 4829 6138 4851
rect 6104 4783 6138 4791
rect 6104 4757 6138 4783
rect 6104 4715 6138 4719
rect 6104 4685 6138 4715
rect 6104 4613 6138 4647
rect 6104 4545 6138 4575
rect 6104 4541 6138 4545
rect 6104 4477 6138 4503
rect 6104 4469 6138 4477
rect 6104 4409 6138 4431
rect 6104 4397 6138 4409
rect 6104 4341 6138 4359
rect 6104 4325 6138 4341
rect 6104 4273 6138 4287
rect 6104 4253 6138 4273
rect 6104 4205 6138 4215
rect 6104 4181 6138 4205
rect 6104 4137 6138 4143
rect 6104 4109 6138 4137
rect 6104 4069 6138 4071
rect 6104 4037 6138 4069
rect 6104 3967 6138 3999
rect 6104 3965 6138 3967
rect 6104 3899 6138 3927
rect 6104 3893 6138 3899
rect 6104 3831 6138 3855
rect 6104 3821 6138 3831
rect 6104 3763 6138 3783
rect 6104 3749 6138 3763
rect 6104 3695 6138 3711
rect 6104 3677 6138 3695
rect 6546 5565 6580 5583
rect 6546 5549 6580 5565
rect 6546 5497 6580 5511
rect 6546 5477 6580 5497
rect 6546 5429 6580 5439
rect 6546 5405 6580 5429
rect 6546 5361 6580 5367
rect 6546 5333 6580 5361
rect 6546 5293 6580 5295
rect 6546 5261 6580 5293
rect 6546 5191 6580 5223
rect 6546 5189 6580 5191
rect 6546 5123 6580 5151
rect 6546 5117 6580 5123
rect 6546 5055 6580 5079
rect 6546 5045 6580 5055
rect 6546 4987 6580 5007
rect 6546 4973 6580 4987
rect 6546 4919 6580 4935
rect 6546 4901 6580 4919
rect 6546 4851 6580 4863
rect 6546 4829 6580 4851
rect 6546 4783 6580 4791
rect 6546 4757 6580 4783
rect 6546 4715 6580 4719
rect 6546 4685 6580 4715
rect 6546 4613 6580 4647
rect 6546 4545 6580 4575
rect 6546 4541 6580 4545
rect 6546 4477 6580 4503
rect 6546 4469 6580 4477
rect 6546 4409 6580 4431
rect 6546 4397 6580 4409
rect 6546 4341 6580 4359
rect 6546 4325 6580 4341
rect 6546 4273 6580 4287
rect 6546 4253 6580 4273
rect 6546 4205 6580 4215
rect 6546 4181 6580 4205
rect 6546 4137 6580 4143
rect 6546 4109 6580 4137
rect 6546 4069 6580 4071
rect 6546 4037 6580 4069
rect 6546 3967 6580 3999
rect 6546 3965 6580 3967
rect 6546 3899 6580 3927
rect 6546 3893 6580 3899
rect 6546 3831 6580 3855
rect 6546 3821 6580 3831
rect 6546 3763 6580 3783
rect 6546 3749 6580 3763
rect 6546 3695 6580 3711
rect 6546 3677 6580 3695
rect 6804 5565 6838 5583
rect 6804 5549 6838 5565
rect 6804 5497 6838 5511
rect 6804 5477 6838 5497
rect 6804 5429 6838 5439
rect 6804 5405 6838 5429
rect 6804 5361 6838 5367
rect 6804 5333 6838 5361
rect 6804 5293 6838 5295
rect 6804 5261 6838 5293
rect 6804 5191 6838 5223
rect 6804 5189 6838 5191
rect 6804 5123 6838 5151
rect 6804 5117 6838 5123
rect 6804 5055 6838 5079
rect 6804 5045 6838 5055
rect 6804 4987 6838 5007
rect 6804 4973 6838 4987
rect 6804 4919 6838 4935
rect 6804 4901 6838 4919
rect 6804 4851 6838 4863
rect 6804 4829 6838 4851
rect 6804 4783 6838 4791
rect 6804 4757 6838 4783
rect 6804 4715 6838 4719
rect 6804 4685 6838 4715
rect 6804 4613 6838 4647
rect 6804 4545 6838 4575
rect 6804 4541 6838 4545
rect 6804 4477 6838 4503
rect 6804 4469 6838 4477
rect 6804 4409 6838 4431
rect 6804 4397 6838 4409
rect 6804 4341 6838 4359
rect 6804 4325 6838 4341
rect 6804 4273 6838 4287
rect 6804 4253 6838 4273
rect 6804 4205 6838 4215
rect 6804 4181 6838 4205
rect 6804 4137 6838 4143
rect 6804 4109 6838 4137
rect 6804 4069 6838 4071
rect 6804 4037 6838 4069
rect 6804 3967 6838 3999
rect 6804 3965 6838 3967
rect 6804 3899 6838 3927
rect 6804 3893 6838 3899
rect 6804 3831 6838 3855
rect 6804 3821 6838 3831
rect 6804 3763 6838 3783
rect 6804 3749 6838 3763
rect 6804 3695 6838 3711
rect 6804 3677 6838 3695
rect 7246 5565 7280 5583
rect 7246 5549 7280 5565
rect 7246 5497 7280 5511
rect 7246 5477 7280 5497
rect 7246 5429 7280 5439
rect 7246 5405 7280 5429
rect 7246 5361 7280 5367
rect 7246 5333 7280 5361
rect 7246 5293 7280 5295
rect 7246 5261 7280 5293
rect 7246 5191 7280 5223
rect 7246 5189 7280 5191
rect 7246 5123 7280 5151
rect 7246 5117 7280 5123
rect 7246 5055 7280 5079
rect 7246 5045 7280 5055
rect 7246 4987 7280 5007
rect 7246 4973 7280 4987
rect 7246 4919 7280 4935
rect 7246 4901 7280 4919
rect 7246 4851 7280 4863
rect 7246 4829 7280 4851
rect 7246 4783 7280 4791
rect 7246 4757 7280 4783
rect 7246 4715 7280 4719
rect 7246 4685 7280 4715
rect 7246 4613 7280 4647
rect 7246 4545 7280 4575
rect 7246 4541 7280 4545
rect 7246 4477 7280 4503
rect 7246 4469 7280 4477
rect 7246 4409 7280 4431
rect 7246 4397 7280 4409
rect 7246 4341 7280 4359
rect 7246 4325 7280 4341
rect 7246 4273 7280 4287
rect 7246 4253 7280 4273
rect 7246 4205 7280 4215
rect 7246 4181 7280 4205
rect 7246 4137 7280 4143
rect 7246 4109 7280 4137
rect 7246 4069 7280 4071
rect 7246 4037 7280 4069
rect 7246 3967 7280 3999
rect 7246 3965 7280 3967
rect 7246 3899 7280 3927
rect 7246 3893 7280 3899
rect 7246 3831 7280 3855
rect 7246 3821 7280 3831
rect 7246 3763 7280 3783
rect 7246 3749 7280 3763
rect 7246 3695 7280 3711
rect 7246 3677 7280 3695
rect 7504 5565 7538 5583
rect 7504 5549 7538 5565
rect 7504 5497 7538 5511
rect 7504 5477 7538 5497
rect 7504 5429 7538 5439
rect 7504 5405 7538 5429
rect 7504 5361 7538 5367
rect 7504 5333 7538 5361
rect 7504 5293 7538 5295
rect 7504 5261 7538 5293
rect 7504 5191 7538 5223
rect 7504 5189 7538 5191
rect 7504 5123 7538 5151
rect 7504 5117 7538 5123
rect 7504 5055 7538 5079
rect 7504 5045 7538 5055
rect 7504 4987 7538 5007
rect 7504 4973 7538 4987
rect 7504 4919 7538 4935
rect 7504 4901 7538 4919
rect 7504 4851 7538 4863
rect 7504 4829 7538 4851
rect 7504 4783 7538 4791
rect 7504 4757 7538 4783
rect 7504 4715 7538 4719
rect 7504 4685 7538 4715
rect 7504 4613 7538 4647
rect 7504 4545 7538 4575
rect 7504 4541 7538 4545
rect 7504 4477 7538 4503
rect 7504 4469 7538 4477
rect 7504 4409 7538 4431
rect 7504 4397 7538 4409
rect 7504 4341 7538 4359
rect 7504 4325 7538 4341
rect 7504 4273 7538 4287
rect 7504 4253 7538 4273
rect 7504 4205 7538 4215
rect 7504 4181 7538 4205
rect 7504 4137 7538 4143
rect 7504 4109 7538 4137
rect 7504 4069 7538 4071
rect 7504 4037 7538 4069
rect 7504 3967 7538 3999
rect 7504 3965 7538 3967
rect 7504 3899 7538 3927
rect 7504 3893 7538 3899
rect 7504 3831 7538 3855
rect 7504 3821 7538 3831
rect 7504 3763 7538 3783
rect 7504 3749 7538 3763
rect 7504 3695 7538 3711
rect 7504 3677 7538 3695
rect 7946 5565 7980 5583
rect 7946 5549 7980 5565
rect 7946 5497 7980 5511
rect 7946 5477 7980 5497
rect 7946 5429 7980 5439
rect 7946 5405 7980 5429
rect 7946 5361 7980 5367
rect 7946 5333 7980 5361
rect 7946 5293 7980 5295
rect 7946 5261 7980 5293
rect 7946 5191 7980 5223
rect 7946 5189 7980 5191
rect 7946 5123 7980 5151
rect 7946 5117 7980 5123
rect 7946 5055 7980 5079
rect 7946 5045 7980 5055
rect 7946 4987 7980 5007
rect 7946 4973 7980 4987
rect 7946 4919 7980 4935
rect 7946 4901 7980 4919
rect 7946 4851 7980 4863
rect 7946 4829 7980 4851
rect 7946 4783 7980 4791
rect 7946 4757 7980 4783
rect 7946 4715 7980 4719
rect 7946 4685 7980 4715
rect 7946 4613 7980 4647
rect 7946 4545 7980 4575
rect 7946 4541 7980 4545
rect 7946 4477 7980 4503
rect 7946 4469 7980 4477
rect 7946 4409 7980 4431
rect 7946 4397 7980 4409
rect 7946 4341 7980 4359
rect 7946 4325 7980 4341
rect 7946 4273 7980 4287
rect 7946 4253 7980 4273
rect 7946 4205 7980 4215
rect 7946 4181 7980 4205
rect 7946 4137 7980 4143
rect 7946 4109 7980 4137
rect 7946 4069 7980 4071
rect 7946 4037 7980 4069
rect 7946 3967 7980 3999
rect 7946 3965 7980 3967
rect 7946 3899 7980 3927
rect 7946 3893 7980 3899
rect 7946 3831 7980 3855
rect 7946 3821 7980 3831
rect 7946 3763 7980 3783
rect 7946 3749 7980 3763
rect 7946 3695 7980 3711
rect 7946 3677 7980 3695
rect 8204 5565 8238 5583
rect 8204 5549 8238 5565
rect 8204 5497 8238 5511
rect 8204 5477 8238 5497
rect 8204 5429 8238 5439
rect 8204 5405 8238 5429
rect 8204 5361 8238 5367
rect 8204 5333 8238 5361
rect 8204 5293 8238 5295
rect 8204 5261 8238 5293
rect 8204 5191 8238 5223
rect 8204 5189 8238 5191
rect 8204 5123 8238 5151
rect 8204 5117 8238 5123
rect 8204 5055 8238 5079
rect 8204 5045 8238 5055
rect 8204 4987 8238 5007
rect 8204 4973 8238 4987
rect 8204 4919 8238 4935
rect 8204 4901 8238 4919
rect 8204 4851 8238 4863
rect 8204 4829 8238 4851
rect 8204 4783 8238 4791
rect 8204 4757 8238 4783
rect 8204 4715 8238 4719
rect 8204 4685 8238 4715
rect 8204 4613 8238 4647
rect 8204 4545 8238 4575
rect 8204 4541 8238 4545
rect 8204 4477 8238 4503
rect 8204 4469 8238 4477
rect 8204 4409 8238 4431
rect 8204 4397 8238 4409
rect 8204 4341 8238 4359
rect 8204 4325 8238 4341
rect 8204 4273 8238 4287
rect 8204 4253 8238 4273
rect 8204 4205 8238 4215
rect 8204 4181 8238 4205
rect 8204 4137 8238 4143
rect 8204 4109 8238 4137
rect 8204 4069 8238 4071
rect 8204 4037 8238 4069
rect 8204 3967 8238 3999
rect 8204 3965 8238 3967
rect 8204 3899 8238 3927
rect 8204 3893 8238 3899
rect 8204 3831 8238 3855
rect 8204 3821 8238 3831
rect 8204 3763 8238 3783
rect 8204 3749 8238 3763
rect 8204 3695 8238 3711
rect 8204 3677 8238 3695
rect 8646 5565 8680 5583
rect 8646 5549 8680 5565
rect 8646 5497 8680 5511
rect 8646 5477 8680 5497
rect 8646 5429 8680 5439
rect 8646 5405 8680 5429
rect 8646 5361 8680 5367
rect 8646 5333 8680 5361
rect 8646 5293 8680 5295
rect 8646 5261 8680 5293
rect 8646 5191 8680 5223
rect 8646 5189 8680 5191
rect 8646 5123 8680 5151
rect 8646 5117 8680 5123
rect 8646 5055 8680 5079
rect 8646 5045 8680 5055
rect 8646 4987 8680 5007
rect 8646 4973 8680 4987
rect 8646 4919 8680 4935
rect 8646 4901 8680 4919
rect 8646 4851 8680 4863
rect 8646 4829 8680 4851
rect 8646 4783 8680 4791
rect 8646 4757 8680 4783
rect 8646 4715 8680 4719
rect 8646 4685 8680 4715
rect 8646 4613 8680 4647
rect 8646 4545 8680 4575
rect 8646 4541 8680 4545
rect 8646 4477 8680 4503
rect 8646 4469 8680 4477
rect 8646 4409 8680 4431
rect 8646 4397 8680 4409
rect 8646 4341 8680 4359
rect 8646 4325 8680 4341
rect 8646 4273 8680 4287
rect 8646 4253 8680 4273
rect 8646 4205 8680 4215
rect 8646 4181 8680 4205
rect 8646 4137 8680 4143
rect 8646 4109 8680 4137
rect 8646 4069 8680 4071
rect 8646 4037 8680 4069
rect 8646 3967 8680 3999
rect 8646 3965 8680 3967
rect 8646 3899 8680 3927
rect 8646 3893 8680 3899
rect 8646 3831 8680 3855
rect 8646 3821 8680 3831
rect 8646 3763 8680 3783
rect 8646 3749 8680 3763
rect 8646 3695 8680 3711
rect 8646 3677 8680 3695
rect 8904 5565 8938 5583
rect 8904 5549 8938 5565
rect 8904 5497 8938 5511
rect 8904 5477 8938 5497
rect 8904 5429 8938 5439
rect 8904 5405 8938 5429
rect 8904 5361 8938 5367
rect 8904 5333 8938 5361
rect 8904 5293 8938 5295
rect 8904 5261 8938 5293
rect 8904 5191 8938 5223
rect 8904 5189 8938 5191
rect 8904 5123 8938 5151
rect 8904 5117 8938 5123
rect 8904 5055 8938 5079
rect 8904 5045 8938 5055
rect 8904 4987 8938 5007
rect 8904 4973 8938 4987
rect 8904 4919 8938 4935
rect 8904 4901 8938 4919
rect 8904 4851 8938 4863
rect 8904 4829 8938 4851
rect 8904 4783 8938 4791
rect 8904 4757 8938 4783
rect 8904 4715 8938 4719
rect 8904 4685 8938 4715
rect 8904 4613 8938 4647
rect 8904 4545 8938 4575
rect 8904 4541 8938 4545
rect 8904 4477 8938 4503
rect 8904 4469 8938 4477
rect 8904 4409 8938 4431
rect 8904 4397 8938 4409
rect 8904 4341 8938 4359
rect 8904 4325 8938 4341
rect 8904 4273 8938 4287
rect 8904 4253 8938 4273
rect 8904 4205 8938 4215
rect 8904 4181 8938 4205
rect 8904 4137 8938 4143
rect 8904 4109 8938 4137
rect 8904 4069 8938 4071
rect 8904 4037 8938 4069
rect 8904 3967 8938 3999
rect 8904 3965 8938 3967
rect 8904 3899 8938 3927
rect 8904 3893 8938 3899
rect 8904 3831 8938 3855
rect 8904 3821 8938 3831
rect 8904 3763 8938 3783
rect 8904 3749 8938 3763
rect 8904 3695 8938 3711
rect 8904 3677 8938 3695
rect 9346 5565 9380 5583
rect 9346 5549 9380 5565
rect 9346 5497 9380 5511
rect 9346 5477 9380 5497
rect 9346 5429 9380 5439
rect 9346 5405 9380 5429
rect 9346 5361 9380 5367
rect 9346 5333 9380 5361
rect 9346 5293 9380 5295
rect 9346 5261 9380 5293
rect 9346 5191 9380 5223
rect 9346 5189 9380 5191
rect 9346 5123 9380 5151
rect 9346 5117 9380 5123
rect 9346 5055 9380 5079
rect 9346 5045 9380 5055
rect 9346 4987 9380 5007
rect 9346 4973 9380 4987
rect 9346 4919 9380 4935
rect 9346 4901 9380 4919
rect 9346 4851 9380 4863
rect 9346 4829 9380 4851
rect 9346 4783 9380 4791
rect 9346 4757 9380 4783
rect 9346 4715 9380 4719
rect 9346 4685 9380 4715
rect 9346 4613 9380 4647
rect 9346 4545 9380 4575
rect 9346 4541 9380 4545
rect 9346 4477 9380 4503
rect 9346 4469 9380 4477
rect 9346 4409 9380 4431
rect 9346 4397 9380 4409
rect 9346 4341 9380 4359
rect 9346 4325 9380 4341
rect 9346 4273 9380 4287
rect 9346 4253 9380 4273
rect 9346 4205 9380 4215
rect 9346 4181 9380 4205
rect 9346 4137 9380 4143
rect 9346 4109 9380 4137
rect 9346 4069 9380 4071
rect 9346 4037 9380 4069
rect 9346 3967 9380 3999
rect 9346 3965 9380 3967
rect 9346 3899 9380 3927
rect 9346 3893 9380 3899
rect 9346 3831 9380 3855
rect 9346 3821 9380 3831
rect 9346 3763 9380 3783
rect 9346 3749 9380 3763
rect 9346 3695 9380 3711
rect 9346 3677 9380 3695
rect 9604 5565 9638 5583
rect 9604 5549 9638 5565
rect 9604 5497 9638 5511
rect 9604 5477 9638 5497
rect 9604 5429 9638 5439
rect 9604 5405 9638 5429
rect 9604 5361 9638 5367
rect 9604 5333 9638 5361
rect 9604 5293 9638 5295
rect 9604 5261 9638 5293
rect 9604 5191 9638 5223
rect 9604 5189 9638 5191
rect 9604 5123 9638 5151
rect 9604 5117 9638 5123
rect 9604 5055 9638 5079
rect 9604 5045 9638 5055
rect 9604 4987 9638 5007
rect 9604 4973 9638 4987
rect 9604 4919 9638 4935
rect 9604 4901 9638 4919
rect 9604 4851 9638 4863
rect 9604 4829 9638 4851
rect 9604 4783 9638 4791
rect 9604 4757 9638 4783
rect 9604 4715 9638 4719
rect 9604 4685 9638 4715
rect 9604 4613 9638 4647
rect 9604 4545 9638 4575
rect 9604 4541 9638 4545
rect 9604 4477 9638 4503
rect 9604 4469 9638 4477
rect 9604 4409 9638 4431
rect 9604 4397 9638 4409
rect 9604 4341 9638 4359
rect 9604 4325 9638 4341
rect 9604 4273 9638 4287
rect 9604 4253 9638 4273
rect 9604 4205 9638 4215
rect 9604 4181 9638 4205
rect 9604 4137 9638 4143
rect 9604 4109 9638 4137
rect 9604 4069 9638 4071
rect 9604 4037 9638 4069
rect 9604 3967 9638 3999
rect 9604 3965 9638 3967
rect 9604 3899 9638 3927
rect 9604 3893 9638 3899
rect 9604 3831 9638 3855
rect 9604 3821 9638 3831
rect 9604 3763 9638 3783
rect 9604 3749 9638 3763
rect 9604 3695 9638 3711
rect 9604 3677 9638 3695
rect 10046 5565 10080 5583
rect 10046 5549 10080 5565
rect 10046 5497 10080 5511
rect 10046 5477 10080 5497
rect 10046 5429 10080 5439
rect 10046 5405 10080 5429
rect 10046 5361 10080 5367
rect 10046 5333 10080 5361
rect 10046 5293 10080 5295
rect 10046 5261 10080 5293
rect 10046 5191 10080 5223
rect 10046 5189 10080 5191
rect 10046 5123 10080 5151
rect 10046 5117 10080 5123
rect 10046 5055 10080 5079
rect 10046 5045 10080 5055
rect 10046 4987 10080 5007
rect 10046 4973 10080 4987
rect 10046 4919 10080 4935
rect 10046 4901 10080 4919
rect 10046 4851 10080 4863
rect 10046 4829 10080 4851
rect 10046 4783 10080 4791
rect 10046 4757 10080 4783
rect 10046 4715 10080 4719
rect 10046 4685 10080 4715
rect 10046 4613 10080 4647
rect 10046 4545 10080 4575
rect 10046 4541 10080 4545
rect 10046 4477 10080 4503
rect 10046 4469 10080 4477
rect 10046 4409 10080 4431
rect 10046 4397 10080 4409
rect 10046 4341 10080 4359
rect 10046 4325 10080 4341
rect 10046 4273 10080 4287
rect 10046 4253 10080 4273
rect 10046 4205 10080 4215
rect 10046 4181 10080 4205
rect 10046 4137 10080 4143
rect 10046 4109 10080 4137
rect 10046 4069 10080 4071
rect 10046 4037 10080 4069
rect 10046 3967 10080 3999
rect 10046 3965 10080 3967
rect 10046 3899 10080 3927
rect 10046 3893 10080 3899
rect 10046 3831 10080 3855
rect 10046 3821 10080 3831
rect 10046 3763 10080 3783
rect 10046 3749 10080 3763
rect 10046 3695 10080 3711
rect 10046 3677 10080 3695
rect 11781 5628 11789 5662
rect 11789 5628 11815 5662
rect 11853 5628 11857 5662
rect 11857 5628 11887 5662
rect 11925 5628 11959 5662
rect 11997 5628 12027 5662
rect 12027 5628 12031 5662
rect 12069 5628 12095 5662
rect 12095 5628 12103 5662
rect 12681 5628 12689 5662
rect 12689 5628 12715 5662
rect 12753 5628 12757 5662
rect 12757 5628 12787 5662
rect 12825 5628 12859 5662
rect 12897 5628 12927 5662
rect 12927 5628 12931 5662
rect 12969 5628 12995 5662
rect 12995 5628 13003 5662
rect 13581 5628 13589 5662
rect 13589 5628 13615 5662
rect 13653 5628 13657 5662
rect 13657 5628 13687 5662
rect 13725 5628 13759 5662
rect 13797 5628 13827 5662
rect 13827 5628 13831 5662
rect 13869 5628 13895 5662
rect 13895 5628 13903 5662
rect 14481 5628 14489 5662
rect 14489 5628 14515 5662
rect 14553 5628 14557 5662
rect 14557 5628 14587 5662
rect 14625 5628 14659 5662
rect 14697 5628 14727 5662
rect 14727 5628 14731 5662
rect 14769 5628 14795 5662
rect 14795 5628 14803 5662
rect 15381 5628 15389 5662
rect 15389 5628 15415 5662
rect 15453 5628 15457 5662
rect 15457 5628 15487 5662
rect 15525 5628 15559 5662
rect 15597 5628 15627 5662
rect 15627 5628 15631 5662
rect 15669 5628 15695 5662
rect 15695 5628 15703 5662
rect 16281 5628 16289 5662
rect 16289 5628 16315 5662
rect 16353 5628 16357 5662
rect 16357 5628 16387 5662
rect 16425 5628 16459 5662
rect 16497 5628 16527 5662
rect 16527 5628 16531 5662
rect 16569 5628 16595 5662
rect 16595 5628 16603 5662
rect 17181 5628 17189 5662
rect 17189 5628 17215 5662
rect 17253 5628 17257 5662
rect 17257 5628 17287 5662
rect 17325 5628 17359 5662
rect 17397 5628 17427 5662
rect 17427 5628 17431 5662
rect 17469 5628 17495 5662
rect 17495 5628 17503 5662
rect 18081 5628 18089 5662
rect 18089 5628 18115 5662
rect 18153 5628 18157 5662
rect 18157 5628 18187 5662
rect 18225 5628 18259 5662
rect 18297 5628 18327 5662
rect 18327 5628 18331 5662
rect 18369 5628 18395 5662
rect 18395 5628 18403 5662
rect 10304 5565 10338 5583
rect 10304 5549 10338 5565
rect 10304 5497 10338 5511
rect 10304 5477 10338 5497
rect 11882 5455 11916 5489
rect 11954 5455 11988 5489
rect 12782 5455 12816 5489
rect 12854 5455 12888 5489
rect 13682 5455 13716 5489
rect 13754 5455 13788 5489
rect 14582 5455 14616 5489
rect 14654 5455 14688 5489
rect 15482 5455 15516 5489
rect 15554 5455 15588 5489
rect 16382 5455 16416 5489
rect 16454 5455 16488 5489
rect 17282 5455 17316 5489
rect 17354 5455 17388 5489
rect 18182 5455 18216 5489
rect 18254 5455 18288 5489
rect 10304 5429 10338 5439
rect 10304 5405 10338 5429
rect 10304 5361 10338 5367
rect 10304 5333 10338 5361
rect 10304 5293 10338 5295
rect 10304 5261 10338 5293
rect 10304 5191 10338 5223
rect 10304 5189 10338 5191
rect 10304 5123 10338 5151
rect 10304 5117 10338 5123
rect 10304 5055 10338 5079
rect 10304 5045 10338 5055
rect 10304 4987 10338 5007
rect 10304 4973 10338 4987
rect 10304 4919 10338 4935
rect 10304 4901 10338 4919
rect 10304 4851 10338 4863
rect 10304 4829 10338 4851
rect 10304 4783 10338 4791
rect 10304 4757 10338 4783
rect 10304 4715 10338 4719
rect 10304 4685 10338 4715
rect 10304 4613 10338 4647
rect 10304 4545 10338 4575
rect 10304 4541 10338 4545
rect 10304 4477 10338 4503
rect 10304 4469 10338 4477
rect 10304 4409 10338 4431
rect 10304 4397 10338 4409
rect 10304 4341 10338 4359
rect 10304 4325 10338 4341
rect 10304 4273 10338 4287
rect 10304 4253 10338 4273
rect 10304 4205 10338 4215
rect 10304 4181 10338 4205
rect 10304 4137 10338 4143
rect 10304 4109 10338 4137
rect 10304 4069 10338 4071
rect 10304 4037 10338 4069
rect 10304 3967 10338 3999
rect 10304 3965 10338 3967
rect 10304 3899 10338 3927
rect 10304 3893 10338 3899
rect 10304 3831 10338 3855
rect 10304 3821 10338 3831
rect 10304 3763 10338 3783
rect 10304 3749 10338 3763
rect 10304 3695 10338 3711
rect 10304 3677 10338 3695
rect -4161 3558 -4159 3592
rect -4159 3558 -4127 3592
rect -4089 3558 -4057 3592
rect -4057 3558 -4055 3592
rect -3461 3558 -3459 3592
rect -3459 3558 -3427 3592
rect -3389 3558 -3357 3592
rect -3357 3558 -3355 3592
rect -2761 3558 -2759 3592
rect -2759 3558 -2727 3592
rect -2689 3558 -2657 3592
rect -2657 3558 -2655 3592
rect -2061 3558 -2059 3592
rect -2059 3558 -2027 3592
rect -1989 3558 -1957 3592
rect -1957 3558 -1955 3592
rect -1361 3558 -1359 3592
rect -1359 3558 -1327 3592
rect -1289 3558 -1257 3592
rect -1257 3558 -1255 3592
rect -661 3558 -659 3592
rect -659 3558 -627 3592
rect -589 3558 -557 3592
rect -557 3558 -555 3592
rect 39 3558 41 3592
rect 41 3558 73 3592
rect 111 3558 143 3592
rect 143 3558 145 3592
rect 739 3558 741 3592
rect 741 3558 773 3592
rect 811 3558 843 3592
rect 843 3558 845 3592
rect 1439 3558 1441 3592
rect 1441 3558 1473 3592
rect 1511 3558 1543 3592
rect 1543 3558 1545 3592
rect 2139 3558 2141 3592
rect 2141 3558 2173 3592
rect 2211 3558 2243 3592
rect 2243 3558 2245 3592
rect 3839 3558 3841 3592
rect 3841 3558 3873 3592
rect 3911 3558 3943 3592
rect 3943 3558 3945 3592
rect 4539 3558 4541 3592
rect 4541 3558 4573 3592
rect 4611 3558 4643 3592
rect 4643 3558 4645 3592
rect 5239 3558 5241 3592
rect 5241 3558 5273 3592
rect 5311 3558 5343 3592
rect 5343 3558 5345 3592
rect 5939 3558 5941 3592
rect 5941 3558 5973 3592
rect 6011 3558 6043 3592
rect 6043 3558 6045 3592
rect 6639 3558 6641 3592
rect 6641 3558 6673 3592
rect 6711 3558 6743 3592
rect 6743 3558 6745 3592
rect 7339 3558 7341 3592
rect 7341 3558 7373 3592
rect 7411 3558 7443 3592
rect 7443 3558 7445 3592
rect 8039 3558 8041 3592
rect 8041 3558 8073 3592
rect 8111 3558 8143 3592
rect 8143 3558 8145 3592
rect 8739 3558 8741 3592
rect 8741 3558 8773 3592
rect 8811 3558 8843 3592
rect 8843 3558 8845 3592
rect 9439 3558 9441 3592
rect 9441 3558 9473 3592
rect 9511 3558 9543 3592
rect 9543 3558 9545 3592
rect 10139 3558 10141 3592
rect 10141 3558 10173 3592
rect 10211 3558 10243 3592
rect 10243 3558 10245 3592
rect 1285 2100 1319 2134
rect 1357 2100 1391 2134
rect 2285 2100 2319 2134
rect 2357 2100 2391 2134
rect 3285 2100 3319 2134
rect 3357 2100 3391 2134
rect 4285 2100 4319 2134
rect 4357 2100 4391 2134
rect 5285 2100 5319 2134
rect 5357 2100 5391 2134
rect 6285 2100 6319 2134
rect 6357 2100 6391 2134
rect 7285 2100 7319 2134
rect 7357 2100 7391 2134
rect 8285 2100 8319 2134
rect 8357 2100 8391 2134
rect 9285 2100 9319 2134
rect 9357 2100 9391 2134
rect 10285 2100 10319 2134
rect 10357 2100 10391 2134
rect 1173 1954 1181 1988
rect 1181 1954 1207 1988
rect 1245 1954 1249 1988
rect 1249 1954 1279 1988
rect 1317 1954 1351 1988
rect 1389 1954 1419 1988
rect 1419 1954 1423 1988
rect 1461 1954 1487 1988
rect 1487 1954 1495 1988
rect 2173 1954 2181 1988
rect 2181 1954 2207 1988
rect 2245 1954 2249 1988
rect 2249 1954 2279 1988
rect 2317 1954 2351 1988
rect 2389 1954 2419 1988
rect 2419 1954 2423 1988
rect 2461 1954 2487 1988
rect 2487 1954 2495 1988
rect 3173 1954 3181 1988
rect 3181 1954 3207 1988
rect 3245 1954 3249 1988
rect 3249 1954 3279 1988
rect 3317 1954 3351 1988
rect 3389 1954 3419 1988
rect 3419 1954 3423 1988
rect 3461 1954 3487 1988
rect 3487 1954 3495 1988
rect 4173 1954 4181 1988
rect 4181 1954 4207 1988
rect 4245 1954 4249 1988
rect 4249 1954 4279 1988
rect 4317 1954 4351 1988
rect 4389 1954 4419 1988
rect 4419 1954 4423 1988
rect 4461 1954 4487 1988
rect 4487 1954 4495 1988
rect 5173 1954 5181 1988
rect 5181 1954 5207 1988
rect 5245 1954 5249 1988
rect 5249 1954 5279 1988
rect 5317 1954 5351 1988
rect 5389 1954 5419 1988
rect 5419 1954 5423 1988
rect 5461 1954 5487 1988
rect 5487 1954 5495 1988
rect 6173 1954 6181 1988
rect 6181 1954 6207 1988
rect 6245 1954 6249 1988
rect 6249 1954 6279 1988
rect 6317 1954 6351 1988
rect 6389 1954 6419 1988
rect 6419 1954 6423 1988
rect 6461 1954 6487 1988
rect 6487 1954 6495 1988
rect 7173 1954 7181 1988
rect 7181 1954 7207 1988
rect 7245 1954 7249 1988
rect 7249 1954 7279 1988
rect 7317 1954 7351 1988
rect 7389 1954 7419 1988
rect 7419 1954 7423 1988
rect 7461 1954 7487 1988
rect 7487 1954 7495 1988
rect 8173 1954 8181 1988
rect 8181 1954 8207 1988
rect 8245 1954 8249 1988
rect 8249 1954 8279 1988
rect 8317 1954 8351 1988
rect 8389 1954 8419 1988
rect 8419 1954 8423 1988
rect 8461 1954 8487 1988
rect 8487 1954 8495 1988
rect 9173 1954 9181 1988
rect 9181 1954 9207 1988
rect 9245 1954 9249 1988
rect 9249 1954 9279 1988
rect 9317 1954 9351 1988
rect 9389 1954 9419 1988
rect 9419 1954 9423 1988
rect 9461 1954 9487 1988
rect 9487 1954 9495 1988
rect 10173 1954 10181 1988
rect 10181 1954 10207 1988
rect 10245 1954 10249 1988
rect 10249 1954 10279 1988
rect 10317 1954 10351 1988
rect 10389 1954 10419 1988
rect 10419 1954 10423 1988
rect 10461 1954 10487 1988
rect 10487 1954 10495 1988
rect 1088 1867 1122 1869
rect 1088 1835 1122 1867
rect 1088 1765 1122 1797
rect 1088 1763 1122 1765
rect 1546 1867 1580 1869
rect 1546 1835 1580 1867
rect 1546 1765 1580 1797
rect 1546 1763 1580 1765
rect 2088 1867 2122 1869
rect 2088 1835 2122 1867
rect 2088 1765 2122 1797
rect 2088 1763 2122 1765
rect 2546 1867 2580 1869
rect 2546 1835 2580 1867
rect 2546 1765 2580 1797
rect 2546 1763 2580 1765
rect 3088 1867 3122 1869
rect 3088 1835 3122 1867
rect 3088 1765 3122 1797
rect 3088 1763 3122 1765
rect 3546 1867 3580 1869
rect 3546 1835 3580 1867
rect 3546 1765 3580 1797
rect 3546 1763 3580 1765
rect 4088 1867 4122 1869
rect 4088 1835 4122 1867
rect 4088 1765 4122 1797
rect 4088 1763 4122 1765
rect 4546 1867 4580 1869
rect 4546 1835 4580 1867
rect 4546 1765 4580 1797
rect 4546 1763 4580 1765
rect 5088 1867 5122 1869
rect 5088 1835 5122 1867
rect 5088 1765 5122 1797
rect 5088 1763 5122 1765
rect 5546 1867 5580 1869
rect 5546 1835 5580 1867
rect 5546 1765 5580 1797
rect 5546 1763 5580 1765
rect 6088 1867 6122 1869
rect 6088 1835 6122 1867
rect 6088 1765 6122 1797
rect 6088 1763 6122 1765
rect 6546 1867 6580 1869
rect 6546 1835 6580 1867
rect 6546 1765 6580 1797
rect 6546 1763 6580 1765
rect 7088 1867 7122 1869
rect 7088 1835 7122 1867
rect 7088 1765 7122 1797
rect 7088 1763 7122 1765
rect 7546 1867 7580 1869
rect 7546 1835 7580 1867
rect 7546 1765 7580 1797
rect 7546 1763 7580 1765
rect 8088 1867 8122 1869
rect 8088 1835 8122 1867
rect 8088 1765 8122 1797
rect 8088 1763 8122 1765
rect 8546 1867 8580 1869
rect 8546 1835 8580 1867
rect 8546 1765 8580 1797
rect 8546 1763 8580 1765
rect 9088 1867 9122 1869
rect 9088 1835 9122 1867
rect 9088 1765 9122 1797
rect 9088 1763 9122 1765
rect 9546 1867 9580 1869
rect 9546 1835 9580 1867
rect 9546 1765 9580 1797
rect 9546 1763 9580 1765
rect 10088 1867 10122 1869
rect 10088 1835 10122 1867
rect 10088 1765 10122 1797
rect 10088 1763 10122 1765
rect 10546 1867 10580 1869
rect 10546 1835 10580 1867
rect 10546 1765 10580 1797
rect 10546 1763 10580 1765
rect 1173 1644 1181 1678
rect 1181 1644 1207 1678
rect 1245 1644 1249 1678
rect 1249 1644 1279 1678
rect 1317 1644 1351 1678
rect 1389 1644 1419 1678
rect 1419 1644 1423 1678
rect 1461 1644 1487 1678
rect 1487 1644 1495 1678
rect 2173 1644 2181 1678
rect 2181 1644 2207 1678
rect 2245 1644 2249 1678
rect 2249 1644 2279 1678
rect 2317 1644 2351 1678
rect 2389 1644 2419 1678
rect 2419 1644 2423 1678
rect 2461 1644 2487 1678
rect 2487 1644 2495 1678
rect 3173 1644 3181 1678
rect 3181 1644 3207 1678
rect 3245 1644 3249 1678
rect 3249 1644 3279 1678
rect 3317 1644 3351 1678
rect 3389 1644 3419 1678
rect 3419 1644 3423 1678
rect 3461 1644 3487 1678
rect 3487 1644 3495 1678
rect 4173 1644 4181 1678
rect 4181 1644 4207 1678
rect 4245 1644 4249 1678
rect 4249 1644 4279 1678
rect 4317 1644 4351 1678
rect 4389 1644 4419 1678
rect 4419 1644 4423 1678
rect 4461 1644 4487 1678
rect 4487 1644 4495 1678
rect 5173 1644 5181 1678
rect 5181 1644 5207 1678
rect 5245 1644 5249 1678
rect 5249 1644 5279 1678
rect 5317 1644 5351 1678
rect 5389 1644 5419 1678
rect 5419 1644 5423 1678
rect 5461 1644 5487 1678
rect 5487 1644 5495 1678
rect 6173 1644 6181 1678
rect 6181 1644 6207 1678
rect 6245 1644 6249 1678
rect 6249 1644 6279 1678
rect 6317 1644 6351 1678
rect 6389 1644 6419 1678
rect 6419 1644 6423 1678
rect 6461 1644 6487 1678
rect 6487 1644 6495 1678
rect 7173 1644 7181 1678
rect 7181 1644 7207 1678
rect 7245 1644 7249 1678
rect 7249 1644 7279 1678
rect 7317 1644 7351 1678
rect 7389 1644 7419 1678
rect 7419 1644 7423 1678
rect 7461 1644 7487 1678
rect 7487 1644 7495 1678
rect 8173 1644 8181 1678
rect 8181 1644 8207 1678
rect 8245 1644 8249 1678
rect 8249 1644 8279 1678
rect 8317 1644 8351 1678
rect 8389 1644 8419 1678
rect 8419 1644 8423 1678
rect 8461 1644 8487 1678
rect 8487 1644 8495 1678
rect 9173 1644 9181 1678
rect 9181 1644 9207 1678
rect 9245 1644 9249 1678
rect 9249 1644 9279 1678
rect 9317 1644 9351 1678
rect 9389 1644 9419 1678
rect 9419 1644 9423 1678
rect 9461 1644 9487 1678
rect 9487 1644 9495 1678
rect 10173 1644 10181 1678
rect 10181 1644 10207 1678
rect 10245 1644 10249 1678
rect 10249 1644 10279 1678
rect 10317 1644 10351 1678
rect 10389 1644 10419 1678
rect 10419 1644 10423 1678
rect 10461 1644 10487 1678
rect 10487 1644 10495 1678
rect 1173 1454 1181 1488
rect 1181 1454 1207 1488
rect 1245 1454 1249 1488
rect 1249 1454 1279 1488
rect 1317 1454 1351 1488
rect 1389 1454 1419 1488
rect 1419 1454 1423 1488
rect 1461 1454 1487 1488
rect 1487 1454 1495 1488
rect 2173 1454 2181 1488
rect 2181 1454 2207 1488
rect 2245 1454 2249 1488
rect 2249 1454 2279 1488
rect 2317 1454 2351 1488
rect 2389 1454 2419 1488
rect 2419 1454 2423 1488
rect 2461 1454 2487 1488
rect 2487 1454 2495 1488
rect 3173 1454 3181 1488
rect 3181 1454 3207 1488
rect 3245 1454 3249 1488
rect 3249 1454 3279 1488
rect 3317 1454 3351 1488
rect 3389 1454 3419 1488
rect 3419 1454 3423 1488
rect 3461 1454 3487 1488
rect 3487 1454 3495 1488
rect 4173 1454 4181 1488
rect 4181 1454 4207 1488
rect 4245 1454 4249 1488
rect 4249 1454 4279 1488
rect 4317 1454 4351 1488
rect 4389 1454 4419 1488
rect 4419 1454 4423 1488
rect 4461 1454 4487 1488
rect 4487 1454 4495 1488
rect 5173 1454 5181 1488
rect 5181 1454 5207 1488
rect 5245 1454 5249 1488
rect 5249 1454 5279 1488
rect 5317 1454 5351 1488
rect 5389 1454 5419 1488
rect 5419 1454 5423 1488
rect 5461 1454 5487 1488
rect 5487 1454 5495 1488
rect 6173 1454 6181 1488
rect 6181 1454 6207 1488
rect 6245 1454 6249 1488
rect 6249 1454 6279 1488
rect 6317 1454 6351 1488
rect 6389 1454 6419 1488
rect 6419 1454 6423 1488
rect 6461 1454 6487 1488
rect 6487 1454 6495 1488
rect 7173 1454 7181 1488
rect 7181 1454 7207 1488
rect 7245 1454 7249 1488
rect 7249 1454 7279 1488
rect 7317 1454 7351 1488
rect 7389 1454 7419 1488
rect 7419 1454 7423 1488
rect 7461 1454 7487 1488
rect 7487 1454 7495 1488
rect 8173 1454 8181 1488
rect 8181 1454 8207 1488
rect 8245 1454 8249 1488
rect 8249 1454 8279 1488
rect 8317 1454 8351 1488
rect 8389 1454 8419 1488
rect 8419 1454 8423 1488
rect 8461 1454 8487 1488
rect 8487 1454 8495 1488
rect 9173 1454 9181 1488
rect 9181 1454 9207 1488
rect 9245 1454 9249 1488
rect 9249 1454 9279 1488
rect 9317 1454 9351 1488
rect 9389 1454 9419 1488
rect 9419 1454 9423 1488
rect 9461 1454 9487 1488
rect 9487 1454 9495 1488
rect 10173 1454 10181 1488
rect 10181 1454 10207 1488
rect 10245 1454 10249 1488
rect 10249 1454 10279 1488
rect 10317 1454 10351 1488
rect 10389 1454 10419 1488
rect 10419 1454 10423 1488
rect 10461 1454 10487 1488
rect 10487 1454 10495 1488
rect 1088 1367 1122 1369
rect 1088 1335 1122 1367
rect 1088 1265 1122 1297
rect 1088 1263 1122 1265
rect 1546 1367 1580 1369
rect 1546 1335 1580 1367
rect 1546 1265 1580 1297
rect 1546 1263 1580 1265
rect 2088 1367 2122 1369
rect 2088 1335 2122 1367
rect 2088 1265 2122 1297
rect 2088 1263 2122 1265
rect 2546 1367 2580 1369
rect 2546 1335 2580 1367
rect 2546 1265 2580 1297
rect 2546 1263 2580 1265
rect 3088 1367 3122 1369
rect 3088 1335 3122 1367
rect 3088 1265 3122 1297
rect 3088 1263 3122 1265
rect 3546 1367 3580 1369
rect 3546 1335 3580 1367
rect 3546 1265 3580 1297
rect 3546 1263 3580 1265
rect 4088 1367 4122 1369
rect 4088 1335 4122 1367
rect 4088 1265 4122 1297
rect 4088 1263 4122 1265
rect 4546 1367 4580 1369
rect 4546 1335 4580 1367
rect 4546 1265 4580 1297
rect 4546 1263 4580 1265
rect 5088 1367 5122 1369
rect 5088 1335 5122 1367
rect 5088 1265 5122 1297
rect 5088 1263 5122 1265
rect 5546 1367 5580 1369
rect 5546 1335 5580 1367
rect 5546 1265 5580 1297
rect 5546 1263 5580 1265
rect 6088 1367 6122 1369
rect 6088 1335 6122 1367
rect 6088 1265 6122 1297
rect 6088 1263 6122 1265
rect 6546 1367 6580 1369
rect 6546 1335 6580 1367
rect 6546 1265 6580 1297
rect 6546 1263 6580 1265
rect 7088 1367 7122 1369
rect 7088 1335 7122 1367
rect 7088 1265 7122 1297
rect 7088 1263 7122 1265
rect 7546 1367 7580 1369
rect 7546 1335 7580 1367
rect 7546 1265 7580 1297
rect 7546 1263 7580 1265
rect 8088 1367 8122 1369
rect 8088 1335 8122 1367
rect 8088 1265 8122 1297
rect 8088 1263 8122 1265
rect 8546 1367 8580 1369
rect 8546 1335 8580 1367
rect 8546 1265 8580 1297
rect 8546 1263 8580 1265
rect 9088 1367 9122 1369
rect 9088 1335 9122 1367
rect 9088 1265 9122 1297
rect 9088 1263 9122 1265
rect 9546 1367 9580 1369
rect 9546 1335 9580 1367
rect 9546 1265 9580 1297
rect 9546 1263 9580 1265
rect 10088 1367 10122 1369
rect 10088 1335 10122 1367
rect 10088 1265 10122 1297
rect 10088 1263 10122 1265
rect 10546 1367 10580 1369
rect 10546 1335 10580 1367
rect 10546 1265 10580 1297
rect 10546 1263 10580 1265
rect 1173 1144 1181 1178
rect 1181 1144 1207 1178
rect 1245 1144 1249 1178
rect 1249 1144 1279 1178
rect 1317 1144 1351 1178
rect 1389 1144 1419 1178
rect 1419 1144 1423 1178
rect 1461 1144 1487 1178
rect 1487 1144 1495 1178
rect 2173 1144 2181 1178
rect 2181 1144 2207 1178
rect 2245 1144 2249 1178
rect 2249 1144 2279 1178
rect 2317 1144 2351 1178
rect 2389 1144 2419 1178
rect 2419 1144 2423 1178
rect 2461 1144 2487 1178
rect 2487 1144 2495 1178
rect 3173 1144 3181 1178
rect 3181 1144 3207 1178
rect 3245 1144 3249 1178
rect 3249 1144 3279 1178
rect 3317 1144 3351 1178
rect 3389 1144 3419 1178
rect 3419 1144 3423 1178
rect 3461 1144 3487 1178
rect 3487 1144 3495 1178
rect 4173 1144 4181 1178
rect 4181 1144 4207 1178
rect 4245 1144 4249 1178
rect 4249 1144 4279 1178
rect 4317 1144 4351 1178
rect 4389 1144 4419 1178
rect 4419 1144 4423 1178
rect 4461 1144 4487 1178
rect 4487 1144 4495 1178
rect 5173 1144 5181 1178
rect 5181 1144 5207 1178
rect 5245 1144 5249 1178
rect 5249 1144 5279 1178
rect 5317 1144 5351 1178
rect 5389 1144 5419 1178
rect 5419 1144 5423 1178
rect 5461 1144 5487 1178
rect 5487 1144 5495 1178
rect 6173 1144 6181 1178
rect 6181 1144 6207 1178
rect 6245 1144 6249 1178
rect 6249 1144 6279 1178
rect 6317 1144 6351 1178
rect 6389 1144 6419 1178
rect 6419 1144 6423 1178
rect 6461 1144 6487 1178
rect 6487 1144 6495 1178
rect 7173 1144 7181 1178
rect 7181 1144 7207 1178
rect 7245 1144 7249 1178
rect 7249 1144 7279 1178
rect 7317 1144 7351 1178
rect 7389 1144 7419 1178
rect 7419 1144 7423 1178
rect 7461 1144 7487 1178
rect 7487 1144 7495 1178
rect 8173 1144 8181 1178
rect 8181 1144 8207 1178
rect 8245 1144 8249 1178
rect 8249 1144 8279 1178
rect 8317 1144 8351 1178
rect 8389 1144 8419 1178
rect 8419 1144 8423 1178
rect 8461 1144 8487 1178
rect 8487 1144 8495 1178
rect 9173 1144 9181 1178
rect 9181 1144 9207 1178
rect 9245 1144 9249 1178
rect 9249 1144 9279 1178
rect 9317 1144 9351 1178
rect 9389 1144 9419 1178
rect 9419 1144 9423 1178
rect 9461 1144 9487 1178
rect 9487 1144 9495 1178
rect 10173 1144 10181 1178
rect 10181 1144 10207 1178
rect 10245 1144 10249 1178
rect 10249 1144 10279 1178
rect 10317 1144 10351 1178
rect 10389 1144 10419 1178
rect 10419 1144 10423 1178
rect 10461 1144 10487 1178
rect 10487 1144 10495 1178
rect 1284 963 1318 997
rect 1356 963 1390 997
rect 2284 963 2318 997
rect 2356 963 2390 997
rect 3284 963 3318 997
rect 3356 963 3390 997
rect 4284 963 4318 997
rect 4356 963 4390 997
rect 5284 963 5318 997
rect 5356 963 5390 997
rect 6284 963 6318 997
rect 6356 963 6390 997
rect 7284 963 7318 997
rect 7356 963 7390 997
rect 8284 963 8318 997
rect 8356 963 8390 997
rect 9284 963 9318 997
rect 9356 963 9390 997
rect 10284 963 10318 997
rect 10356 963 10390 997
<< metal1 >>
rect -9200 8951 4266 9070
rect -9200 8950 -9080 8951
rect 1839 8789 1972 8951
rect 2839 8789 2972 8951
rect 1839 8754 2300 8789
rect 1839 8720 2167 8754
rect 2201 8720 2239 8754
rect 2273 8720 2300 8754
rect 1839 8685 2300 8720
rect 2839 8754 3300 8789
rect 2839 8720 3167 8754
rect 3201 8720 3239 8754
rect 3273 8720 3300 8754
rect 2839 8685 3300 8720
rect 1839 8509 1972 8685
rect 2028 8590 2420 8596
rect 2028 8556 2063 8590
rect 2097 8556 2135 8590
rect 2169 8556 2207 8590
rect 2241 8556 2279 8590
rect 2313 8556 2351 8590
rect 2385 8556 2420 8590
rect 2028 8550 2420 8556
rect 2476 8509 2609 8640
rect 1839 8470 2018 8509
rect 1839 8436 1978 8470
rect 2012 8436 2018 8470
rect 1839 8398 2018 8436
rect 1839 8364 1978 8398
rect 2012 8364 2018 8398
rect 1839 8326 2018 8364
rect 1839 8292 1978 8326
rect 2012 8292 2018 8326
rect 1839 8254 2018 8292
rect 1839 8220 1978 8254
rect 2012 8220 2018 8254
rect 1839 8182 2018 8220
rect 1839 8148 1978 8182
rect 2012 8148 2018 8182
rect 1839 8109 2018 8148
rect 2430 8470 2609 8509
rect 2430 8436 2436 8470
rect 2470 8436 2609 8470
rect 2430 8398 2609 8436
rect 2430 8364 2436 8398
rect 2470 8364 2609 8398
rect 2430 8326 2609 8364
rect 2430 8292 2436 8326
rect 2470 8292 2609 8326
rect 2430 8254 2609 8292
rect 2430 8220 2436 8254
rect 2470 8220 2609 8254
rect 2430 8182 2609 8220
rect 2430 8148 2436 8182
rect 2470 8148 2609 8182
rect 2430 8109 2609 8148
rect 1839 7769 1972 8109
rect 2028 8062 2420 8068
rect 2028 8028 2063 8062
rect 2097 8028 2135 8062
rect 2169 8028 2207 8062
rect 2241 8028 2279 8062
rect 2313 8028 2351 8062
rect 2385 8028 2420 8062
rect 2028 8022 2420 8028
rect 2476 8022 2609 8109
rect 2028 7969 2609 8022
rect 2028 7917 2176 7969
rect 2228 7917 2240 7969
rect 2292 7917 2609 7969
rect 2028 7856 2609 7917
rect 2028 7850 2420 7856
rect 2028 7816 2063 7850
rect 2097 7816 2135 7850
rect 2169 7816 2207 7850
rect 2241 7816 2279 7850
rect 2313 7816 2351 7850
rect 2385 7816 2420 7850
rect 2028 7810 2420 7816
rect 2476 7769 2609 7856
rect 1839 7730 2018 7769
rect 1839 7696 1978 7730
rect 2012 7696 2018 7730
rect 1839 7658 2018 7696
rect 1839 7624 1978 7658
rect 2012 7624 2018 7658
rect 1839 7586 2018 7624
rect 1839 7552 1978 7586
rect 2012 7552 2018 7586
rect 1839 7514 2018 7552
rect 1839 7480 1978 7514
rect 2012 7480 2018 7514
rect 1839 7442 2018 7480
rect 1839 7408 1978 7442
rect 2012 7408 2018 7442
rect 1839 7369 2018 7408
rect 2430 7730 2609 7769
rect 2430 7696 2436 7730
rect 2470 7696 2609 7730
rect 2430 7658 2609 7696
rect 2430 7624 2436 7658
rect 2470 7624 2609 7658
rect 2430 7586 2609 7624
rect 2430 7552 2436 7586
rect 2470 7552 2609 7586
rect 2430 7514 2609 7552
rect 2430 7480 2436 7514
rect 2470 7480 2609 7514
rect 2430 7442 2609 7480
rect 2430 7408 2436 7442
rect 2470 7408 2609 7442
rect 2430 7369 2609 7408
rect 1839 7184 1972 7369
rect 2028 7322 2420 7328
rect 2028 7288 2063 7322
rect 2097 7288 2135 7322
rect 2169 7288 2207 7322
rect 2241 7288 2279 7322
rect 2313 7288 2351 7322
rect 2385 7288 2420 7322
rect 2028 7282 2420 7288
rect 1839 7149 2300 7184
rect 1839 7115 2164 7149
rect 2198 7115 2236 7149
rect 2270 7115 2300 7149
rect 1839 7080 2300 7115
rect 2476 6413 2609 7369
rect 2839 8509 2972 8685
rect 3028 8590 3420 8596
rect 3028 8556 3063 8590
rect 3097 8556 3135 8590
rect 3169 8556 3207 8590
rect 3241 8556 3279 8590
rect 3313 8556 3351 8590
rect 3385 8556 3420 8590
rect 3028 8550 3420 8556
rect 3476 8509 3609 8640
rect 2839 8470 3018 8509
rect 2839 8436 2978 8470
rect 3012 8436 3018 8470
rect 2839 8398 3018 8436
rect 2839 8364 2978 8398
rect 3012 8364 3018 8398
rect 2839 8326 3018 8364
rect 2839 8292 2978 8326
rect 3012 8292 3018 8326
rect 2839 8254 3018 8292
rect 2839 8220 2978 8254
rect 3012 8220 3018 8254
rect 2839 8182 3018 8220
rect 2839 8148 2978 8182
rect 3012 8148 3018 8182
rect 2839 8109 3018 8148
rect 3430 8470 3609 8509
rect 3430 8436 3436 8470
rect 3470 8436 3609 8470
rect 3430 8398 3609 8436
rect 3430 8364 3436 8398
rect 3470 8364 3609 8398
rect 3430 8326 3609 8364
rect 3430 8292 3436 8326
rect 3470 8292 3609 8326
rect 3430 8254 3609 8292
rect 3430 8220 3436 8254
rect 3470 8220 3609 8254
rect 3430 8182 3609 8220
rect 3430 8148 3436 8182
rect 3470 8148 3609 8182
rect 3430 8109 3609 8148
rect 2839 7769 2972 8109
rect 3028 8062 3420 8068
rect 3028 8028 3063 8062
rect 3097 8028 3135 8062
rect 3169 8028 3207 8062
rect 3241 8028 3279 8062
rect 3313 8028 3351 8062
rect 3385 8028 3420 8062
rect 3028 7969 3420 8028
rect 3028 7917 3176 7969
rect 3228 7917 3240 7969
rect 3292 7917 3420 7969
rect 3028 7850 3420 7917
rect 3028 7816 3063 7850
rect 3097 7816 3135 7850
rect 3169 7816 3207 7850
rect 3241 7816 3279 7850
rect 3313 7816 3351 7850
rect 3385 7816 3420 7850
rect 3028 7810 3420 7816
rect 3476 7769 3609 8109
rect 2839 7730 3018 7769
rect 2839 7696 2978 7730
rect 3012 7696 3018 7730
rect 2839 7658 3018 7696
rect 2839 7624 2978 7658
rect 3012 7624 3018 7658
rect 2839 7586 3018 7624
rect 2839 7552 2978 7586
rect 3012 7552 3018 7586
rect 2839 7514 3018 7552
rect 2839 7480 2978 7514
rect 3012 7480 3018 7514
rect 2839 7442 3018 7480
rect 2839 7408 2978 7442
rect 3012 7408 3018 7442
rect 2839 7369 3018 7408
rect 3430 7730 3609 7769
rect 3430 7696 3436 7730
rect 3470 7696 3609 7730
rect 3430 7658 3609 7696
rect 3430 7624 3436 7658
rect 3470 7624 3609 7658
rect 3430 7586 3609 7624
rect 3430 7552 3436 7586
rect 3470 7552 3609 7586
rect 3430 7514 3609 7552
rect 3430 7480 3436 7514
rect 3470 7480 3609 7514
rect 3430 7442 3609 7480
rect 3430 7408 3436 7442
rect 3470 7408 3609 7442
rect 3430 7369 3609 7408
rect 2839 7184 2972 7369
rect 3028 7322 3420 7328
rect 3028 7288 3063 7322
rect 3097 7288 3135 7322
rect 3169 7288 3207 7322
rect 3241 7288 3279 7322
rect 3313 7288 3351 7322
rect 3385 7288 3420 7322
rect 3028 7282 3420 7288
rect 2839 7149 3300 7184
rect 2839 7115 3164 7149
rect 3198 7115 3236 7149
rect 3270 7115 3300 7149
rect 2839 7080 3300 7115
rect 2012 6340 2614 6413
rect 3476 6409 3609 7369
rect 4125 7474 4266 8951
rect 21449 8900 21567 8914
rect 21449 8506 21455 8900
rect 21561 8506 21567 8900
rect 21449 8493 21567 8506
rect 21073 7602 21155 7627
rect 21073 7568 21097 7602
rect 21131 7568 21155 7602
rect 21073 7530 21155 7568
rect 21073 7496 21097 7530
rect 21131 7496 21155 7530
rect 4125 7291 17990 7474
rect -4396 6182 2614 6340
rect 3477 6340 3609 6409
rect 11557 7129 11690 7291
rect 12457 7129 12590 7291
rect 13357 7129 13490 7291
rect 14257 7129 14390 7291
rect 15157 7129 15290 7291
rect 16057 7129 16190 7291
rect 16957 7129 17090 7291
rect 17857 7129 17990 7291
rect 11557 7094 12018 7129
rect 11557 7060 11885 7094
rect 11919 7060 11957 7094
rect 11991 7060 12018 7094
rect 11557 7025 12018 7060
rect 12457 7094 12918 7129
rect 12457 7060 12785 7094
rect 12819 7060 12857 7094
rect 12891 7060 12918 7094
rect 12457 7025 12918 7060
rect 13357 7094 13818 7129
rect 13357 7060 13685 7094
rect 13719 7060 13757 7094
rect 13791 7060 13818 7094
rect 13357 7025 13818 7060
rect 14257 7094 14718 7129
rect 14257 7060 14585 7094
rect 14619 7060 14657 7094
rect 14691 7060 14718 7094
rect 14257 7025 14718 7060
rect 15157 7094 15618 7129
rect 15157 7060 15485 7094
rect 15519 7060 15557 7094
rect 15591 7060 15618 7094
rect 15157 7025 15618 7060
rect 16057 7094 16518 7129
rect 16057 7060 16385 7094
rect 16419 7060 16457 7094
rect 16491 7060 16518 7094
rect 16057 7025 16518 7060
rect 16957 7094 17418 7129
rect 16957 7060 17285 7094
rect 17319 7060 17357 7094
rect 17391 7060 17418 7094
rect 16957 7025 17418 7060
rect 17857 7094 18318 7129
rect 17857 7060 18185 7094
rect 18219 7060 18257 7094
rect 18291 7060 18318 7094
rect 17857 7025 18318 7060
rect 11557 6849 11690 7025
rect 11746 6930 12138 6936
rect 11746 6896 11781 6930
rect 11815 6896 11853 6930
rect 11887 6896 11925 6930
rect 11959 6896 11997 6930
rect 12031 6896 12069 6930
rect 12103 6896 12138 6930
rect 11746 6890 12138 6896
rect 12194 6849 12327 6980
rect 11557 6810 11736 6849
rect 11557 6776 11696 6810
rect 11730 6776 11736 6810
rect 11557 6738 11736 6776
rect 11557 6704 11696 6738
rect 11730 6704 11736 6738
rect 11557 6666 11736 6704
rect 11557 6632 11696 6666
rect 11730 6632 11736 6666
rect 11557 6594 11736 6632
rect 11557 6560 11696 6594
rect 11730 6560 11736 6594
rect 11557 6522 11736 6560
rect 11557 6488 11696 6522
rect 11730 6488 11736 6522
rect 11557 6449 11736 6488
rect 12148 6810 12327 6849
rect 12148 6776 12154 6810
rect 12188 6776 12327 6810
rect 12148 6738 12327 6776
rect 12148 6704 12154 6738
rect 12188 6704 12327 6738
rect 12148 6666 12327 6704
rect 12148 6632 12154 6666
rect 12188 6632 12327 6666
rect 12148 6594 12327 6632
rect 12148 6560 12154 6594
rect 12188 6560 12327 6594
rect 12148 6522 12327 6560
rect 12148 6488 12154 6522
rect 12188 6488 12327 6522
rect 12148 6449 12327 6488
rect 3477 6310 10040 6340
rect 3477 6304 10060 6310
rect 3477 6252 9938 6304
rect 9990 6252 10002 6304
rect 10054 6252 10060 6304
rect 3477 6246 10060 6252
rect 3477 6188 10040 6246
rect -4396 6180 2040 6182
rect -4794 5942 -4689 5953
rect -4794 5890 -4768 5942
rect -4716 5890 -4689 5942
rect -4794 5878 -4689 5890
rect -4794 5826 -4768 5878
rect -4716 5826 -4689 5878
rect -4794 2751 -4689 5826
rect -4396 5630 -4260 6180
rect -4204 5702 -4012 5708
rect -4204 5668 -4161 5702
rect -4127 5668 -4089 5702
rect -4055 5668 -4012 5702
rect -4204 5662 -4012 5668
rect -3696 5630 -3560 6180
rect -3504 5702 -3312 5708
rect -3504 5668 -3461 5702
rect -3427 5668 -3389 5702
rect -3355 5668 -3312 5702
rect -3504 5662 -3312 5668
rect -2996 5630 -2860 6180
rect -2804 5702 -2612 5708
rect -2804 5668 -2761 5702
rect -2727 5668 -2689 5702
rect -2655 5668 -2612 5702
rect -2804 5662 -2612 5668
rect -2296 5630 -2160 6180
rect -2104 5702 -1912 5708
rect -2104 5668 -2061 5702
rect -2027 5668 -1989 5702
rect -1955 5668 -1912 5702
rect -2104 5662 -1912 5668
rect -1596 5630 -1460 6180
rect -1404 5702 -1212 5708
rect -1404 5668 -1361 5702
rect -1327 5668 -1289 5702
rect -1255 5668 -1212 5702
rect -1404 5662 -1212 5668
rect -896 5630 -760 6180
rect -704 5702 -512 5708
rect -704 5668 -661 5702
rect -627 5668 -589 5702
rect -555 5668 -512 5702
rect -704 5662 -512 5668
rect -196 5630 -60 6180
rect -4 5702 188 5708
rect -4 5668 39 5702
rect 73 5668 111 5702
rect 145 5668 188 5702
rect -4 5662 188 5668
rect 504 5630 640 6180
rect 696 5702 888 5708
rect 696 5668 739 5702
rect 773 5668 811 5702
rect 845 5668 888 5702
rect 696 5662 888 5668
rect 1204 5630 1340 6180
rect 1396 5702 1588 5708
rect 1396 5668 1439 5702
rect 1473 5668 1511 5702
rect 1545 5668 1588 5702
rect 1396 5662 1588 5668
rect 1904 5630 2040 6180
rect 3604 6180 10040 6188
rect 2096 5702 2288 5708
rect 2096 5668 2139 5702
rect 2173 5668 2211 5702
rect 2245 5668 2288 5702
rect 2096 5662 2288 5668
rect 3604 5630 3740 6180
rect 3796 5702 3988 5708
rect 3796 5668 3839 5702
rect 3873 5668 3911 5702
rect 3945 5668 3988 5702
rect 3796 5662 3988 5668
rect 4304 5630 4440 6180
rect 4496 5702 4688 5708
rect 4496 5668 4539 5702
rect 4573 5668 4611 5702
rect 4645 5668 4688 5702
rect 4496 5662 4688 5668
rect 5004 5630 5140 6180
rect 5196 5702 5388 5708
rect 5196 5668 5239 5702
rect 5273 5668 5311 5702
rect 5345 5668 5388 5702
rect 5196 5662 5388 5668
rect 5704 5630 5840 6180
rect 5896 5702 6088 5708
rect 5896 5668 5939 5702
rect 5973 5668 6011 5702
rect 6045 5668 6088 5702
rect 5896 5662 6088 5668
rect 6404 5630 6540 6180
rect 6596 5702 6788 5708
rect 6596 5668 6639 5702
rect 6673 5668 6711 5702
rect 6745 5668 6788 5702
rect 6596 5662 6788 5668
rect 7104 5630 7240 6180
rect 7296 5702 7488 5708
rect 7296 5668 7339 5702
rect 7373 5668 7411 5702
rect 7445 5668 7488 5702
rect 7296 5662 7488 5668
rect 7804 5630 7940 6180
rect 7996 5702 8188 5708
rect 7996 5668 8039 5702
rect 8073 5668 8111 5702
rect 8145 5668 8188 5702
rect 7996 5662 8188 5668
rect 8504 5630 8640 6180
rect 8696 5702 8888 5708
rect 8696 5668 8739 5702
rect 8773 5668 8811 5702
rect 8845 5668 8888 5702
rect 8696 5662 8888 5668
rect 9204 5630 9340 6180
rect 9396 5702 9588 5708
rect 9396 5668 9439 5702
rect 9473 5668 9511 5702
rect 9545 5668 9588 5702
rect 9396 5662 9588 5668
rect 9904 5630 10040 6180
rect 11557 6109 11690 6449
rect 11746 6402 12138 6408
rect 11746 6368 11781 6402
rect 11815 6368 11853 6402
rect 11887 6368 11925 6402
rect 11959 6368 11997 6402
rect 12031 6368 12069 6402
rect 12103 6368 12138 6402
rect 11746 6305 12138 6368
rect 11746 6253 11894 6305
rect 11946 6253 11958 6305
rect 12010 6253 12138 6305
rect 11746 6190 12138 6253
rect 11746 6156 11781 6190
rect 11815 6156 11853 6190
rect 11887 6156 11925 6190
rect 11959 6156 11997 6190
rect 12031 6156 12069 6190
rect 12103 6156 12138 6190
rect 11746 6150 12138 6156
rect 12194 6109 12327 6449
rect 11557 6070 11736 6109
rect 11557 6036 11696 6070
rect 11730 6036 11736 6070
rect 11557 5998 11736 6036
rect 11557 5964 11696 5998
rect 11730 5964 11736 5998
rect 11557 5926 11736 5964
rect 11557 5892 11696 5926
rect 11730 5892 11736 5926
rect 11557 5854 11736 5892
rect 11557 5820 11696 5854
rect 11730 5820 11736 5854
rect 11557 5782 11736 5820
rect 11557 5748 11696 5782
rect 11730 5748 11736 5782
rect 11557 5709 11736 5748
rect 12148 6070 12327 6109
rect 12148 6036 12154 6070
rect 12188 6036 12327 6070
rect 12148 5998 12327 6036
rect 12148 5964 12154 5998
rect 12188 5964 12327 5998
rect 12148 5926 12327 5964
rect 12148 5892 12154 5926
rect 12188 5892 12327 5926
rect 12148 5854 12327 5892
rect 12148 5820 12154 5854
rect 12188 5820 12327 5854
rect 12148 5782 12327 5820
rect 12148 5748 12154 5782
rect 12188 5748 12327 5782
rect 12148 5709 12327 5748
rect 10096 5702 10288 5708
rect 10096 5668 10139 5702
rect 10173 5668 10211 5702
rect 10245 5668 10288 5702
rect 10096 5662 10288 5668
rect -4396 5583 -4214 5630
rect -4396 5549 -4254 5583
rect -4220 5549 -4214 5583
rect -4396 5511 -4214 5549
rect -4396 5477 -4254 5511
rect -4220 5477 -4214 5511
rect -4396 5439 -4214 5477
rect -4396 5405 -4254 5439
rect -4220 5405 -4214 5439
rect -4396 5367 -4214 5405
rect -4396 5333 -4254 5367
rect -4220 5333 -4214 5367
rect -4396 5295 -4214 5333
rect -4396 5261 -4254 5295
rect -4220 5261 -4214 5295
rect -4396 5223 -4214 5261
rect -4396 5189 -4254 5223
rect -4220 5189 -4214 5223
rect -4396 5151 -4214 5189
rect -4396 5117 -4254 5151
rect -4220 5117 -4214 5151
rect -4396 5079 -4214 5117
rect -4396 5045 -4254 5079
rect -4220 5045 -4214 5079
rect -4396 5007 -4214 5045
rect -4396 4973 -4254 5007
rect -4220 4973 -4214 5007
rect -4396 4935 -4214 4973
rect -4396 4901 -4254 4935
rect -4220 4901 -4214 4935
rect -4396 4863 -4214 4901
rect -4396 4829 -4254 4863
rect -4220 4829 -4214 4863
rect -4396 4791 -4214 4829
rect -4396 4757 -4254 4791
rect -4220 4757 -4214 4791
rect -4396 4719 -4214 4757
rect -4396 4685 -4254 4719
rect -4220 4685 -4214 4719
rect -4396 4647 -4214 4685
rect -4396 4613 -4254 4647
rect -4220 4613 -4214 4647
rect -4396 4575 -4214 4613
rect -4396 4541 -4254 4575
rect -4220 4541 -4214 4575
rect -4396 4503 -4214 4541
rect -4396 4469 -4254 4503
rect -4220 4469 -4214 4503
rect -4396 4431 -4214 4469
rect -4396 4397 -4254 4431
rect -4220 4397 -4214 4431
rect -4396 4359 -4214 4397
rect -4396 4325 -4254 4359
rect -4220 4325 -4214 4359
rect -4396 4287 -4214 4325
rect -4396 4253 -4254 4287
rect -4220 4253 -4214 4287
rect -4396 4215 -4214 4253
rect -4396 4181 -4254 4215
rect -4220 4181 -4214 4215
rect -4396 4143 -4214 4181
rect -4396 4109 -4254 4143
rect -4220 4109 -4214 4143
rect -4396 4071 -4214 4109
rect -4396 4037 -4254 4071
rect -4220 4037 -4214 4071
rect -4396 3999 -4214 4037
rect -4396 3965 -4254 3999
rect -4220 3965 -4214 3999
rect -4396 3927 -4214 3965
rect -4396 3893 -4254 3927
rect -4220 3893 -4214 3927
rect -4396 3855 -4214 3893
rect -4396 3821 -4254 3855
rect -4220 3821 -4214 3855
rect -4396 3783 -4214 3821
rect -4396 3749 -4254 3783
rect -4220 3749 -4214 3783
rect -4396 3711 -4214 3749
rect -4396 3677 -4254 3711
rect -4220 3677 -4214 3711
rect -4396 3630 -4214 3677
rect -4002 5583 -3820 5630
rect -4002 5549 -3996 5583
rect -3962 5549 -3820 5583
rect -4002 5511 -3820 5549
rect -4002 5477 -3996 5511
rect -3962 5477 -3820 5511
rect -4002 5439 -3820 5477
rect -4002 5405 -3996 5439
rect -3962 5405 -3820 5439
rect -4002 5367 -3820 5405
rect -4002 5333 -3996 5367
rect -3962 5333 -3820 5367
rect -4002 5295 -3820 5333
rect -4002 5261 -3996 5295
rect -3962 5261 -3820 5295
rect -4002 5223 -3820 5261
rect -4002 5189 -3996 5223
rect -3962 5189 -3820 5223
rect -4002 5151 -3820 5189
rect -4002 5117 -3996 5151
rect -3962 5117 -3820 5151
rect -4002 5079 -3820 5117
rect -4002 5045 -3996 5079
rect -3962 5045 -3820 5079
rect -4002 5007 -3820 5045
rect -4002 4973 -3996 5007
rect -3962 4973 -3820 5007
rect -4002 4935 -3820 4973
rect -4002 4901 -3996 4935
rect -3962 4901 -3820 4935
rect -4002 4863 -3820 4901
rect -4002 4829 -3996 4863
rect -3962 4829 -3820 4863
rect -4002 4791 -3820 4829
rect -4002 4757 -3996 4791
rect -3962 4757 -3820 4791
rect -4002 4719 -3820 4757
rect -4002 4685 -3996 4719
rect -3962 4685 -3820 4719
rect -4002 4647 -3820 4685
rect -4002 4613 -3996 4647
rect -3962 4613 -3820 4647
rect -4002 4575 -3820 4613
rect -4002 4541 -3996 4575
rect -3962 4541 -3820 4575
rect -4002 4503 -3820 4541
rect -4002 4469 -3996 4503
rect -3962 4469 -3820 4503
rect -4002 4431 -3820 4469
rect -4002 4397 -3996 4431
rect -3962 4397 -3820 4431
rect -4002 4359 -3820 4397
rect -4002 4325 -3996 4359
rect -3962 4325 -3820 4359
rect -4002 4287 -3820 4325
rect -4002 4253 -3996 4287
rect -3962 4253 -3820 4287
rect -4002 4215 -3820 4253
rect -4002 4181 -3996 4215
rect -3962 4181 -3820 4215
rect -4002 4143 -3820 4181
rect -4002 4109 -3996 4143
rect -3962 4109 -3820 4143
rect -4002 4071 -3820 4109
rect -4002 4037 -3996 4071
rect -3962 4037 -3820 4071
rect -4002 3999 -3820 4037
rect -4002 3965 -3996 3999
rect -3962 3965 -3820 3999
rect -4002 3927 -3820 3965
rect -4002 3893 -3996 3927
rect -3962 3893 -3820 3927
rect -4002 3855 -3820 3893
rect -4002 3821 -3996 3855
rect -3962 3821 -3820 3855
rect -4002 3783 -3820 3821
rect -4002 3749 -3996 3783
rect -3962 3749 -3820 3783
rect -4002 3711 -3820 3749
rect -4002 3677 -3996 3711
rect -3962 3677 -3820 3711
rect -4002 3630 -3820 3677
rect -3696 5583 -3514 5630
rect -3696 5549 -3554 5583
rect -3520 5549 -3514 5583
rect -3696 5511 -3514 5549
rect -3696 5477 -3554 5511
rect -3520 5477 -3514 5511
rect -3696 5439 -3514 5477
rect -3696 5405 -3554 5439
rect -3520 5405 -3514 5439
rect -3696 5367 -3514 5405
rect -3696 5333 -3554 5367
rect -3520 5333 -3514 5367
rect -3696 5295 -3514 5333
rect -3696 5261 -3554 5295
rect -3520 5261 -3514 5295
rect -3696 5223 -3514 5261
rect -3696 5189 -3554 5223
rect -3520 5189 -3514 5223
rect -3696 5151 -3514 5189
rect -3696 5117 -3554 5151
rect -3520 5117 -3514 5151
rect -3696 5079 -3514 5117
rect -3696 5045 -3554 5079
rect -3520 5045 -3514 5079
rect -3696 5007 -3514 5045
rect -3696 4973 -3554 5007
rect -3520 4973 -3514 5007
rect -3696 4935 -3514 4973
rect -3696 4901 -3554 4935
rect -3520 4901 -3514 4935
rect -3696 4863 -3514 4901
rect -3696 4829 -3554 4863
rect -3520 4829 -3514 4863
rect -3696 4791 -3514 4829
rect -3696 4757 -3554 4791
rect -3520 4757 -3514 4791
rect -3696 4719 -3514 4757
rect -3696 4685 -3554 4719
rect -3520 4685 -3514 4719
rect -3696 4647 -3514 4685
rect -3696 4613 -3554 4647
rect -3520 4613 -3514 4647
rect -3696 4575 -3514 4613
rect -3696 4541 -3554 4575
rect -3520 4541 -3514 4575
rect -3696 4503 -3514 4541
rect -3696 4469 -3554 4503
rect -3520 4469 -3514 4503
rect -3696 4431 -3514 4469
rect -3696 4397 -3554 4431
rect -3520 4397 -3514 4431
rect -3696 4359 -3514 4397
rect -3696 4325 -3554 4359
rect -3520 4325 -3514 4359
rect -3696 4287 -3514 4325
rect -3696 4253 -3554 4287
rect -3520 4253 -3514 4287
rect -3696 4215 -3514 4253
rect -3696 4181 -3554 4215
rect -3520 4181 -3514 4215
rect -3696 4143 -3514 4181
rect -3696 4109 -3554 4143
rect -3520 4109 -3514 4143
rect -3696 4071 -3514 4109
rect -3696 4037 -3554 4071
rect -3520 4037 -3514 4071
rect -3696 3999 -3514 4037
rect -3696 3965 -3554 3999
rect -3520 3965 -3514 3999
rect -3696 3927 -3514 3965
rect -3696 3893 -3554 3927
rect -3520 3893 -3514 3927
rect -3696 3855 -3514 3893
rect -3696 3821 -3554 3855
rect -3520 3821 -3514 3855
rect -3696 3783 -3514 3821
rect -3696 3749 -3554 3783
rect -3520 3749 -3514 3783
rect -3696 3711 -3514 3749
rect -3696 3677 -3554 3711
rect -3520 3677 -3514 3711
rect -3696 3630 -3514 3677
rect -3302 5583 -3120 5630
rect -3302 5549 -3296 5583
rect -3262 5549 -3120 5583
rect -3302 5511 -3120 5549
rect -3302 5477 -3296 5511
rect -3262 5477 -3120 5511
rect -3302 5439 -3120 5477
rect -3302 5405 -3296 5439
rect -3262 5405 -3120 5439
rect -3302 5367 -3120 5405
rect -3302 5333 -3296 5367
rect -3262 5333 -3120 5367
rect -3302 5295 -3120 5333
rect -3302 5261 -3296 5295
rect -3262 5261 -3120 5295
rect -3302 5223 -3120 5261
rect -3302 5189 -3296 5223
rect -3262 5189 -3120 5223
rect -3302 5151 -3120 5189
rect -3302 5117 -3296 5151
rect -3262 5117 -3120 5151
rect -3302 5079 -3120 5117
rect -3302 5045 -3296 5079
rect -3262 5045 -3120 5079
rect -3302 5007 -3120 5045
rect -3302 4973 -3296 5007
rect -3262 4973 -3120 5007
rect -3302 4935 -3120 4973
rect -3302 4901 -3296 4935
rect -3262 4901 -3120 4935
rect -3302 4863 -3120 4901
rect -3302 4829 -3296 4863
rect -3262 4829 -3120 4863
rect -3302 4791 -3120 4829
rect -3302 4757 -3296 4791
rect -3262 4757 -3120 4791
rect -3302 4719 -3120 4757
rect -3302 4685 -3296 4719
rect -3262 4685 -3120 4719
rect -3302 4647 -3120 4685
rect -3302 4613 -3296 4647
rect -3262 4613 -3120 4647
rect -3302 4575 -3120 4613
rect -3302 4541 -3296 4575
rect -3262 4541 -3120 4575
rect -3302 4503 -3120 4541
rect -3302 4469 -3296 4503
rect -3262 4469 -3120 4503
rect -3302 4431 -3120 4469
rect -3302 4397 -3296 4431
rect -3262 4397 -3120 4431
rect -3302 4359 -3120 4397
rect -3302 4325 -3296 4359
rect -3262 4325 -3120 4359
rect -3302 4287 -3120 4325
rect -3302 4253 -3296 4287
rect -3262 4253 -3120 4287
rect -3302 4215 -3120 4253
rect -3302 4181 -3296 4215
rect -3262 4181 -3120 4215
rect -3302 4143 -3120 4181
rect -3302 4109 -3296 4143
rect -3262 4109 -3120 4143
rect -3302 4071 -3120 4109
rect -3302 4037 -3296 4071
rect -3262 4037 -3120 4071
rect -3302 3999 -3120 4037
rect -3302 3965 -3296 3999
rect -3262 3965 -3120 3999
rect -3302 3927 -3120 3965
rect -3302 3893 -3296 3927
rect -3262 3893 -3120 3927
rect -3302 3855 -3120 3893
rect -3302 3821 -3296 3855
rect -3262 3821 -3120 3855
rect -3302 3783 -3120 3821
rect -3302 3749 -3296 3783
rect -3262 3749 -3120 3783
rect -3302 3711 -3120 3749
rect -3302 3677 -3296 3711
rect -3262 3677 -3120 3711
rect -3302 3630 -3120 3677
rect -2996 5583 -2814 5630
rect -2996 5549 -2854 5583
rect -2820 5549 -2814 5583
rect -2996 5511 -2814 5549
rect -2996 5477 -2854 5511
rect -2820 5477 -2814 5511
rect -2996 5439 -2814 5477
rect -2996 5405 -2854 5439
rect -2820 5405 -2814 5439
rect -2996 5367 -2814 5405
rect -2996 5333 -2854 5367
rect -2820 5333 -2814 5367
rect -2996 5295 -2814 5333
rect -2996 5261 -2854 5295
rect -2820 5261 -2814 5295
rect -2996 5223 -2814 5261
rect -2996 5189 -2854 5223
rect -2820 5189 -2814 5223
rect -2996 5151 -2814 5189
rect -2996 5117 -2854 5151
rect -2820 5117 -2814 5151
rect -2996 5079 -2814 5117
rect -2996 5045 -2854 5079
rect -2820 5045 -2814 5079
rect -2996 5007 -2814 5045
rect -2996 4973 -2854 5007
rect -2820 4973 -2814 5007
rect -2996 4935 -2814 4973
rect -2996 4901 -2854 4935
rect -2820 4901 -2814 4935
rect -2996 4863 -2814 4901
rect -2996 4829 -2854 4863
rect -2820 4829 -2814 4863
rect -2996 4791 -2814 4829
rect -2996 4757 -2854 4791
rect -2820 4757 -2814 4791
rect -2996 4719 -2814 4757
rect -2996 4685 -2854 4719
rect -2820 4685 -2814 4719
rect -2996 4647 -2814 4685
rect -2996 4613 -2854 4647
rect -2820 4613 -2814 4647
rect -2996 4575 -2814 4613
rect -2996 4541 -2854 4575
rect -2820 4541 -2814 4575
rect -2996 4503 -2814 4541
rect -2996 4469 -2854 4503
rect -2820 4469 -2814 4503
rect -2996 4431 -2814 4469
rect -2996 4397 -2854 4431
rect -2820 4397 -2814 4431
rect -2996 4359 -2814 4397
rect -2996 4325 -2854 4359
rect -2820 4325 -2814 4359
rect -2996 4287 -2814 4325
rect -2996 4253 -2854 4287
rect -2820 4253 -2814 4287
rect -2996 4215 -2814 4253
rect -2996 4181 -2854 4215
rect -2820 4181 -2814 4215
rect -2996 4143 -2814 4181
rect -2996 4109 -2854 4143
rect -2820 4109 -2814 4143
rect -2996 4071 -2814 4109
rect -2996 4037 -2854 4071
rect -2820 4037 -2814 4071
rect -2996 3999 -2814 4037
rect -2996 3965 -2854 3999
rect -2820 3965 -2814 3999
rect -2996 3927 -2814 3965
rect -2996 3893 -2854 3927
rect -2820 3893 -2814 3927
rect -2996 3855 -2814 3893
rect -2996 3821 -2854 3855
rect -2820 3821 -2814 3855
rect -2996 3783 -2814 3821
rect -2996 3749 -2854 3783
rect -2820 3749 -2814 3783
rect -2996 3711 -2814 3749
rect -2996 3677 -2854 3711
rect -2820 3677 -2814 3711
rect -2996 3630 -2814 3677
rect -2602 5583 -2420 5630
rect -2602 5549 -2596 5583
rect -2562 5549 -2420 5583
rect -2602 5511 -2420 5549
rect -2602 5477 -2596 5511
rect -2562 5477 -2420 5511
rect -2602 5439 -2420 5477
rect -2602 5405 -2596 5439
rect -2562 5405 -2420 5439
rect -2602 5367 -2420 5405
rect -2602 5333 -2596 5367
rect -2562 5333 -2420 5367
rect -2602 5295 -2420 5333
rect -2602 5261 -2596 5295
rect -2562 5261 -2420 5295
rect -2602 5223 -2420 5261
rect -2602 5189 -2596 5223
rect -2562 5189 -2420 5223
rect -2602 5151 -2420 5189
rect -2602 5117 -2596 5151
rect -2562 5117 -2420 5151
rect -2602 5079 -2420 5117
rect -2602 5045 -2596 5079
rect -2562 5045 -2420 5079
rect -2602 5007 -2420 5045
rect -2602 4973 -2596 5007
rect -2562 4973 -2420 5007
rect -2602 4935 -2420 4973
rect -2602 4901 -2596 4935
rect -2562 4901 -2420 4935
rect -2602 4863 -2420 4901
rect -2602 4829 -2596 4863
rect -2562 4829 -2420 4863
rect -2602 4791 -2420 4829
rect -2602 4757 -2596 4791
rect -2562 4757 -2420 4791
rect -2602 4719 -2420 4757
rect -2602 4685 -2596 4719
rect -2562 4685 -2420 4719
rect -2602 4647 -2420 4685
rect -2602 4613 -2596 4647
rect -2562 4613 -2420 4647
rect -2602 4575 -2420 4613
rect -2602 4541 -2596 4575
rect -2562 4541 -2420 4575
rect -2602 4503 -2420 4541
rect -2602 4469 -2596 4503
rect -2562 4469 -2420 4503
rect -2602 4431 -2420 4469
rect -2602 4397 -2596 4431
rect -2562 4397 -2420 4431
rect -2602 4359 -2420 4397
rect -2602 4325 -2596 4359
rect -2562 4325 -2420 4359
rect -2602 4287 -2420 4325
rect -2602 4253 -2596 4287
rect -2562 4253 -2420 4287
rect -2602 4215 -2420 4253
rect -2602 4181 -2596 4215
rect -2562 4181 -2420 4215
rect -2602 4143 -2420 4181
rect -2602 4109 -2596 4143
rect -2562 4109 -2420 4143
rect -2602 4071 -2420 4109
rect -2602 4037 -2596 4071
rect -2562 4037 -2420 4071
rect -2602 3999 -2420 4037
rect -2602 3965 -2596 3999
rect -2562 3965 -2420 3999
rect -2602 3927 -2420 3965
rect -2602 3893 -2596 3927
rect -2562 3893 -2420 3927
rect -2602 3855 -2420 3893
rect -2602 3821 -2596 3855
rect -2562 3821 -2420 3855
rect -2602 3783 -2420 3821
rect -2602 3749 -2596 3783
rect -2562 3749 -2420 3783
rect -2602 3711 -2420 3749
rect -2602 3677 -2596 3711
rect -2562 3677 -2420 3711
rect -2602 3630 -2420 3677
rect -2296 5583 -2114 5630
rect -2296 5549 -2154 5583
rect -2120 5549 -2114 5583
rect -2296 5511 -2114 5549
rect -2296 5477 -2154 5511
rect -2120 5477 -2114 5511
rect -2296 5439 -2114 5477
rect -2296 5405 -2154 5439
rect -2120 5405 -2114 5439
rect -2296 5367 -2114 5405
rect -2296 5333 -2154 5367
rect -2120 5333 -2114 5367
rect -2296 5295 -2114 5333
rect -2296 5261 -2154 5295
rect -2120 5261 -2114 5295
rect -2296 5223 -2114 5261
rect -2296 5189 -2154 5223
rect -2120 5189 -2114 5223
rect -2296 5151 -2114 5189
rect -2296 5117 -2154 5151
rect -2120 5117 -2114 5151
rect -2296 5079 -2114 5117
rect -2296 5045 -2154 5079
rect -2120 5045 -2114 5079
rect -2296 5007 -2114 5045
rect -2296 4973 -2154 5007
rect -2120 4973 -2114 5007
rect -2296 4935 -2114 4973
rect -2296 4901 -2154 4935
rect -2120 4901 -2114 4935
rect -2296 4863 -2114 4901
rect -2296 4829 -2154 4863
rect -2120 4829 -2114 4863
rect -2296 4791 -2114 4829
rect -2296 4757 -2154 4791
rect -2120 4757 -2114 4791
rect -2296 4719 -2114 4757
rect -2296 4685 -2154 4719
rect -2120 4685 -2114 4719
rect -2296 4647 -2114 4685
rect -2296 4613 -2154 4647
rect -2120 4613 -2114 4647
rect -2296 4575 -2114 4613
rect -2296 4541 -2154 4575
rect -2120 4541 -2114 4575
rect -2296 4503 -2114 4541
rect -2296 4469 -2154 4503
rect -2120 4469 -2114 4503
rect -2296 4431 -2114 4469
rect -2296 4397 -2154 4431
rect -2120 4397 -2114 4431
rect -2296 4359 -2114 4397
rect -2296 4325 -2154 4359
rect -2120 4325 -2114 4359
rect -2296 4287 -2114 4325
rect -2296 4253 -2154 4287
rect -2120 4253 -2114 4287
rect -2296 4215 -2114 4253
rect -2296 4181 -2154 4215
rect -2120 4181 -2114 4215
rect -2296 4143 -2114 4181
rect -2296 4109 -2154 4143
rect -2120 4109 -2114 4143
rect -2296 4071 -2114 4109
rect -2296 4037 -2154 4071
rect -2120 4037 -2114 4071
rect -2296 3999 -2114 4037
rect -2296 3965 -2154 3999
rect -2120 3965 -2114 3999
rect -2296 3927 -2114 3965
rect -2296 3893 -2154 3927
rect -2120 3893 -2114 3927
rect -2296 3855 -2114 3893
rect -2296 3821 -2154 3855
rect -2120 3821 -2114 3855
rect -2296 3783 -2114 3821
rect -2296 3749 -2154 3783
rect -2120 3749 -2114 3783
rect -2296 3711 -2114 3749
rect -2296 3677 -2154 3711
rect -2120 3677 -2114 3711
rect -2296 3630 -2114 3677
rect -1902 5583 -1720 5630
rect -1902 5549 -1896 5583
rect -1862 5549 -1720 5583
rect -1902 5511 -1720 5549
rect -1902 5477 -1896 5511
rect -1862 5477 -1720 5511
rect -1902 5439 -1720 5477
rect -1902 5405 -1896 5439
rect -1862 5405 -1720 5439
rect -1902 5367 -1720 5405
rect -1902 5333 -1896 5367
rect -1862 5333 -1720 5367
rect -1902 5295 -1720 5333
rect -1902 5261 -1896 5295
rect -1862 5261 -1720 5295
rect -1902 5223 -1720 5261
rect -1902 5189 -1896 5223
rect -1862 5189 -1720 5223
rect -1902 5151 -1720 5189
rect -1902 5117 -1896 5151
rect -1862 5117 -1720 5151
rect -1902 5079 -1720 5117
rect -1902 5045 -1896 5079
rect -1862 5045 -1720 5079
rect -1902 5007 -1720 5045
rect -1902 4973 -1896 5007
rect -1862 4973 -1720 5007
rect -1902 4935 -1720 4973
rect -1902 4901 -1896 4935
rect -1862 4901 -1720 4935
rect -1902 4863 -1720 4901
rect -1902 4829 -1896 4863
rect -1862 4829 -1720 4863
rect -1902 4791 -1720 4829
rect -1902 4757 -1896 4791
rect -1862 4757 -1720 4791
rect -1902 4719 -1720 4757
rect -1902 4685 -1896 4719
rect -1862 4685 -1720 4719
rect -1902 4647 -1720 4685
rect -1902 4613 -1896 4647
rect -1862 4613 -1720 4647
rect -1902 4575 -1720 4613
rect -1902 4541 -1896 4575
rect -1862 4541 -1720 4575
rect -1902 4503 -1720 4541
rect -1902 4469 -1896 4503
rect -1862 4469 -1720 4503
rect -1902 4431 -1720 4469
rect -1902 4397 -1896 4431
rect -1862 4397 -1720 4431
rect -1902 4359 -1720 4397
rect -1902 4325 -1896 4359
rect -1862 4325 -1720 4359
rect -1902 4287 -1720 4325
rect -1902 4253 -1896 4287
rect -1862 4253 -1720 4287
rect -1902 4215 -1720 4253
rect -1902 4181 -1896 4215
rect -1862 4181 -1720 4215
rect -1902 4143 -1720 4181
rect -1902 4109 -1896 4143
rect -1862 4109 -1720 4143
rect -1902 4071 -1720 4109
rect -1902 4037 -1896 4071
rect -1862 4037 -1720 4071
rect -1902 3999 -1720 4037
rect -1902 3965 -1896 3999
rect -1862 3965 -1720 3999
rect -1902 3927 -1720 3965
rect -1902 3893 -1896 3927
rect -1862 3893 -1720 3927
rect -1902 3855 -1720 3893
rect -1902 3821 -1896 3855
rect -1862 3821 -1720 3855
rect -1902 3783 -1720 3821
rect -1902 3749 -1896 3783
rect -1862 3749 -1720 3783
rect -1902 3711 -1720 3749
rect -1902 3677 -1896 3711
rect -1862 3677 -1720 3711
rect -1902 3630 -1720 3677
rect -1596 5583 -1414 5630
rect -1596 5549 -1454 5583
rect -1420 5549 -1414 5583
rect -1596 5511 -1414 5549
rect -1596 5477 -1454 5511
rect -1420 5477 -1414 5511
rect -1596 5439 -1414 5477
rect -1596 5405 -1454 5439
rect -1420 5405 -1414 5439
rect -1596 5367 -1414 5405
rect -1596 5333 -1454 5367
rect -1420 5333 -1414 5367
rect -1596 5295 -1414 5333
rect -1596 5261 -1454 5295
rect -1420 5261 -1414 5295
rect -1596 5223 -1414 5261
rect -1596 5189 -1454 5223
rect -1420 5189 -1414 5223
rect -1596 5151 -1414 5189
rect -1596 5117 -1454 5151
rect -1420 5117 -1414 5151
rect -1596 5079 -1414 5117
rect -1596 5045 -1454 5079
rect -1420 5045 -1414 5079
rect -1596 5007 -1414 5045
rect -1596 4973 -1454 5007
rect -1420 4973 -1414 5007
rect -1596 4935 -1414 4973
rect -1596 4901 -1454 4935
rect -1420 4901 -1414 4935
rect -1596 4863 -1414 4901
rect -1596 4829 -1454 4863
rect -1420 4829 -1414 4863
rect -1596 4791 -1414 4829
rect -1596 4757 -1454 4791
rect -1420 4757 -1414 4791
rect -1596 4719 -1414 4757
rect -1596 4685 -1454 4719
rect -1420 4685 -1414 4719
rect -1596 4647 -1414 4685
rect -1596 4613 -1454 4647
rect -1420 4613 -1414 4647
rect -1596 4575 -1414 4613
rect -1596 4541 -1454 4575
rect -1420 4541 -1414 4575
rect -1596 4503 -1414 4541
rect -1596 4469 -1454 4503
rect -1420 4469 -1414 4503
rect -1596 4431 -1414 4469
rect -1596 4397 -1454 4431
rect -1420 4397 -1414 4431
rect -1596 4359 -1414 4397
rect -1596 4325 -1454 4359
rect -1420 4325 -1414 4359
rect -1596 4287 -1414 4325
rect -1596 4253 -1454 4287
rect -1420 4253 -1414 4287
rect -1596 4215 -1414 4253
rect -1596 4181 -1454 4215
rect -1420 4181 -1414 4215
rect -1596 4143 -1414 4181
rect -1596 4109 -1454 4143
rect -1420 4109 -1414 4143
rect -1596 4071 -1414 4109
rect -1596 4037 -1454 4071
rect -1420 4037 -1414 4071
rect -1596 3999 -1414 4037
rect -1596 3965 -1454 3999
rect -1420 3965 -1414 3999
rect -1596 3927 -1414 3965
rect -1596 3893 -1454 3927
rect -1420 3893 -1414 3927
rect -1596 3855 -1414 3893
rect -1596 3821 -1454 3855
rect -1420 3821 -1414 3855
rect -1596 3783 -1414 3821
rect -1596 3749 -1454 3783
rect -1420 3749 -1414 3783
rect -1596 3711 -1414 3749
rect -1596 3677 -1454 3711
rect -1420 3677 -1414 3711
rect -1596 3630 -1414 3677
rect -1202 5583 -1020 5630
rect -1202 5549 -1196 5583
rect -1162 5549 -1020 5583
rect -1202 5511 -1020 5549
rect -1202 5477 -1196 5511
rect -1162 5477 -1020 5511
rect -1202 5439 -1020 5477
rect -1202 5405 -1196 5439
rect -1162 5405 -1020 5439
rect -1202 5367 -1020 5405
rect -1202 5333 -1196 5367
rect -1162 5333 -1020 5367
rect -1202 5295 -1020 5333
rect -1202 5261 -1196 5295
rect -1162 5261 -1020 5295
rect -1202 5223 -1020 5261
rect -1202 5189 -1196 5223
rect -1162 5189 -1020 5223
rect -1202 5151 -1020 5189
rect -1202 5117 -1196 5151
rect -1162 5117 -1020 5151
rect -1202 5079 -1020 5117
rect -1202 5045 -1196 5079
rect -1162 5045 -1020 5079
rect -1202 5007 -1020 5045
rect -1202 4973 -1196 5007
rect -1162 4973 -1020 5007
rect -1202 4935 -1020 4973
rect -1202 4901 -1196 4935
rect -1162 4901 -1020 4935
rect -1202 4863 -1020 4901
rect -1202 4829 -1196 4863
rect -1162 4829 -1020 4863
rect -1202 4791 -1020 4829
rect -1202 4757 -1196 4791
rect -1162 4757 -1020 4791
rect -1202 4719 -1020 4757
rect -1202 4685 -1196 4719
rect -1162 4685 -1020 4719
rect -1202 4647 -1020 4685
rect -1202 4613 -1196 4647
rect -1162 4613 -1020 4647
rect -1202 4575 -1020 4613
rect -1202 4541 -1196 4575
rect -1162 4541 -1020 4575
rect -1202 4503 -1020 4541
rect -1202 4469 -1196 4503
rect -1162 4469 -1020 4503
rect -1202 4431 -1020 4469
rect -1202 4397 -1196 4431
rect -1162 4397 -1020 4431
rect -1202 4359 -1020 4397
rect -1202 4325 -1196 4359
rect -1162 4325 -1020 4359
rect -1202 4287 -1020 4325
rect -1202 4253 -1196 4287
rect -1162 4253 -1020 4287
rect -1202 4215 -1020 4253
rect -1202 4181 -1196 4215
rect -1162 4181 -1020 4215
rect -1202 4143 -1020 4181
rect -1202 4109 -1196 4143
rect -1162 4109 -1020 4143
rect -1202 4071 -1020 4109
rect -1202 4037 -1196 4071
rect -1162 4037 -1020 4071
rect -1202 3999 -1020 4037
rect -1202 3965 -1196 3999
rect -1162 3965 -1020 3999
rect -1202 3927 -1020 3965
rect -1202 3893 -1196 3927
rect -1162 3893 -1020 3927
rect -1202 3855 -1020 3893
rect -1202 3821 -1196 3855
rect -1162 3821 -1020 3855
rect -1202 3783 -1020 3821
rect -1202 3749 -1196 3783
rect -1162 3749 -1020 3783
rect -1202 3711 -1020 3749
rect -1202 3677 -1196 3711
rect -1162 3677 -1020 3711
rect -1202 3630 -1020 3677
rect -896 5583 -714 5630
rect -896 5549 -754 5583
rect -720 5549 -714 5583
rect -896 5511 -714 5549
rect -896 5477 -754 5511
rect -720 5477 -714 5511
rect -896 5439 -714 5477
rect -896 5405 -754 5439
rect -720 5405 -714 5439
rect -896 5367 -714 5405
rect -896 5333 -754 5367
rect -720 5333 -714 5367
rect -896 5295 -714 5333
rect -896 5261 -754 5295
rect -720 5261 -714 5295
rect -896 5223 -714 5261
rect -896 5189 -754 5223
rect -720 5189 -714 5223
rect -896 5151 -714 5189
rect -896 5117 -754 5151
rect -720 5117 -714 5151
rect -896 5079 -714 5117
rect -896 5045 -754 5079
rect -720 5045 -714 5079
rect -896 5007 -714 5045
rect -896 4973 -754 5007
rect -720 4973 -714 5007
rect -896 4935 -714 4973
rect -896 4901 -754 4935
rect -720 4901 -714 4935
rect -896 4863 -714 4901
rect -896 4829 -754 4863
rect -720 4829 -714 4863
rect -896 4791 -714 4829
rect -896 4757 -754 4791
rect -720 4757 -714 4791
rect -896 4719 -714 4757
rect -896 4685 -754 4719
rect -720 4685 -714 4719
rect -896 4647 -714 4685
rect -896 4613 -754 4647
rect -720 4613 -714 4647
rect -896 4575 -714 4613
rect -896 4541 -754 4575
rect -720 4541 -714 4575
rect -896 4503 -714 4541
rect -896 4469 -754 4503
rect -720 4469 -714 4503
rect -896 4431 -714 4469
rect -896 4397 -754 4431
rect -720 4397 -714 4431
rect -896 4359 -714 4397
rect -896 4325 -754 4359
rect -720 4325 -714 4359
rect -896 4287 -714 4325
rect -896 4253 -754 4287
rect -720 4253 -714 4287
rect -896 4215 -714 4253
rect -896 4181 -754 4215
rect -720 4181 -714 4215
rect -896 4143 -714 4181
rect -896 4109 -754 4143
rect -720 4109 -714 4143
rect -896 4071 -714 4109
rect -896 4037 -754 4071
rect -720 4037 -714 4071
rect -896 3999 -714 4037
rect -896 3965 -754 3999
rect -720 3965 -714 3999
rect -896 3927 -714 3965
rect -896 3893 -754 3927
rect -720 3893 -714 3927
rect -896 3855 -714 3893
rect -896 3821 -754 3855
rect -720 3821 -714 3855
rect -896 3783 -714 3821
rect -896 3749 -754 3783
rect -720 3749 -714 3783
rect -896 3711 -714 3749
rect -896 3677 -754 3711
rect -720 3677 -714 3711
rect -896 3630 -714 3677
rect -502 5583 -320 5630
rect -502 5549 -496 5583
rect -462 5549 -320 5583
rect -502 5511 -320 5549
rect -502 5477 -496 5511
rect -462 5477 -320 5511
rect -502 5439 -320 5477
rect -502 5405 -496 5439
rect -462 5405 -320 5439
rect -502 5367 -320 5405
rect -502 5333 -496 5367
rect -462 5333 -320 5367
rect -502 5295 -320 5333
rect -502 5261 -496 5295
rect -462 5261 -320 5295
rect -502 5223 -320 5261
rect -502 5189 -496 5223
rect -462 5189 -320 5223
rect -502 5151 -320 5189
rect -502 5117 -496 5151
rect -462 5117 -320 5151
rect -502 5079 -320 5117
rect -502 5045 -496 5079
rect -462 5045 -320 5079
rect -502 5007 -320 5045
rect -502 4973 -496 5007
rect -462 4973 -320 5007
rect -502 4935 -320 4973
rect -502 4901 -496 4935
rect -462 4901 -320 4935
rect -502 4863 -320 4901
rect -502 4829 -496 4863
rect -462 4829 -320 4863
rect -502 4791 -320 4829
rect -502 4757 -496 4791
rect -462 4757 -320 4791
rect -502 4719 -320 4757
rect -502 4685 -496 4719
rect -462 4685 -320 4719
rect -502 4647 -320 4685
rect -502 4613 -496 4647
rect -462 4613 -320 4647
rect -502 4575 -320 4613
rect -502 4541 -496 4575
rect -462 4541 -320 4575
rect -502 4503 -320 4541
rect -502 4469 -496 4503
rect -462 4469 -320 4503
rect -502 4431 -320 4469
rect -502 4397 -496 4431
rect -462 4397 -320 4431
rect -502 4359 -320 4397
rect -502 4325 -496 4359
rect -462 4325 -320 4359
rect -502 4287 -320 4325
rect -502 4253 -496 4287
rect -462 4253 -320 4287
rect -502 4215 -320 4253
rect -502 4181 -496 4215
rect -462 4181 -320 4215
rect -502 4143 -320 4181
rect -502 4109 -496 4143
rect -462 4109 -320 4143
rect -502 4071 -320 4109
rect -502 4037 -496 4071
rect -462 4037 -320 4071
rect -502 3999 -320 4037
rect -502 3965 -496 3999
rect -462 3965 -320 3999
rect -502 3927 -320 3965
rect -502 3893 -496 3927
rect -462 3893 -320 3927
rect -502 3855 -320 3893
rect -502 3821 -496 3855
rect -462 3821 -320 3855
rect -502 3783 -320 3821
rect -502 3749 -496 3783
rect -462 3749 -320 3783
rect -502 3711 -320 3749
rect -502 3677 -496 3711
rect -462 3677 -320 3711
rect -502 3630 -320 3677
rect -196 5583 -14 5630
rect -196 5549 -54 5583
rect -20 5549 -14 5583
rect -196 5511 -14 5549
rect -196 5477 -54 5511
rect -20 5477 -14 5511
rect -196 5439 -14 5477
rect -196 5405 -54 5439
rect -20 5405 -14 5439
rect -196 5367 -14 5405
rect -196 5333 -54 5367
rect -20 5333 -14 5367
rect -196 5295 -14 5333
rect -196 5261 -54 5295
rect -20 5261 -14 5295
rect -196 5223 -14 5261
rect -196 5189 -54 5223
rect -20 5189 -14 5223
rect -196 5151 -14 5189
rect -196 5117 -54 5151
rect -20 5117 -14 5151
rect -196 5079 -14 5117
rect -196 5045 -54 5079
rect -20 5045 -14 5079
rect -196 5007 -14 5045
rect -196 4973 -54 5007
rect -20 4973 -14 5007
rect -196 4935 -14 4973
rect -196 4901 -54 4935
rect -20 4901 -14 4935
rect -196 4863 -14 4901
rect -196 4829 -54 4863
rect -20 4829 -14 4863
rect -196 4791 -14 4829
rect -196 4757 -54 4791
rect -20 4757 -14 4791
rect -196 4719 -14 4757
rect -196 4685 -54 4719
rect -20 4685 -14 4719
rect -196 4647 -14 4685
rect -196 4613 -54 4647
rect -20 4613 -14 4647
rect -196 4575 -14 4613
rect -196 4541 -54 4575
rect -20 4541 -14 4575
rect -196 4503 -14 4541
rect -196 4469 -54 4503
rect -20 4469 -14 4503
rect -196 4431 -14 4469
rect -196 4397 -54 4431
rect -20 4397 -14 4431
rect -196 4359 -14 4397
rect -196 4325 -54 4359
rect -20 4325 -14 4359
rect -196 4287 -14 4325
rect -196 4253 -54 4287
rect -20 4253 -14 4287
rect -196 4215 -14 4253
rect -196 4181 -54 4215
rect -20 4181 -14 4215
rect -196 4143 -14 4181
rect -196 4109 -54 4143
rect -20 4109 -14 4143
rect -196 4071 -14 4109
rect -196 4037 -54 4071
rect -20 4037 -14 4071
rect -196 3999 -14 4037
rect -196 3965 -54 3999
rect -20 3965 -14 3999
rect -196 3927 -14 3965
rect -196 3893 -54 3927
rect -20 3893 -14 3927
rect -196 3855 -14 3893
rect -196 3821 -54 3855
rect -20 3821 -14 3855
rect -196 3783 -14 3821
rect -196 3749 -54 3783
rect -20 3749 -14 3783
rect -196 3711 -14 3749
rect -196 3677 -54 3711
rect -20 3677 -14 3711
rect -196 3630 -14 3677
rect 198 5583 380 5630
rect 198 5549 204 5583
rect 238 5549 380 5583
rect 198 5511 380 5549
rect 198 5477 204 5511
rect 238 5477 380 5511
rect 198 5439 380 5477
rect 198 5405 204 5439
rect 238 5405 380 5439
rect 198 5367 380 5405
rect 198 5333 204 5367
rect 238 5333 380 5367
rect 198 5295 380 5333
rect 198 5261 204 5295
rect 238 5261 380 5295
rect 198 5223 380 5261
rect 198 5189 204 5223
rect 238 5189 380 5223
rect 198 5151 380 5189
rect 198 5117 204 5151
rect 238 5117 380 5151
rect 198 5079 380 5117
rect 198 5045 204 5079
rect 238 5045 380 5079
rect 198 5007 380 5045
rect 198 4973 204 5007
rect 238 4973 380 5007
rect 198 4935 380 4973
rect 198 4901 204 4935
rect 238 4901 380 4935
rect 198 4863 380 4901
rect 198 4829 204 4863
rect 238 4829 380 4863
rect 198 4791 380 4829
rect 198 4757 204 4791
rect 238 4757 380 4791
rect 198 4719 380 4757
rect 198 4685 204 4719
rect 238 4685 380 4719
rect 198 4647 380 4685
rect 198 4613 204 4647
rect 238 4613 380 4647
rect 198 4575 380 4613
rect 198 4541 204 4575
rect 238 4541 380 4575
rect 198 4503 380 4541
rect 198 4469 204 4503
rect 238 4469 380 4503
rect 198 4431 380 4469
rect 198 4397 204 4431
rect 238 4397 380 4431
rect 198 4359 380 4397
rect 198 4325 204 4359
rect 238 4325 380 4359
rect 198 4287 380 4325
rect 198 4253 204 4287
rect 238 4253 380 4287
rect 198 4215 380 4253
rect 198 4181 204 4215
rect 238 4181 380 4215
rect 198 4143 380 4181
rect 198 4109 204 4143
rect 238 4109 380 4143
rect 198 4071 380 4109
rect 198 4037 204 4071
rect 238 4037 380 4071
rect 198 3999 380 4037
rect 198 3965 204 3999
rect 238 3965 380 3999
rect 198 3927 380 3965
rect 198 3893 204 3927
rect 238 3893 380 3927
rect 198 3855 380 3893
rect 198 3821 204 3855
rect 238 3821 380 3855
rect 198 3783 380 3821
rect 198 3749 204 3783
rect 238 3749 380 3783
rect 198 3711 380 3749
rect 198 3677 204 3711
rect 238 3677 380 3711
rect 198 3630 380 3677
rect 504 5583 686 5630
rect 504 5549 646 5583
rect 680 5549 686 5583
rect 504 5511 686 5549
rect 504 5477 646 5511
rect 680 5477 686 5511
rect 504 5439 686 5477
rect 504 5405 646 5439
rect 680 5405 686 5439
rect 504 5367 686 5405
rect 504 5333 646 5367
rect 680 5333 686 5367
rect 504 5295 686 5333
rect 504 5261 646 5295
rect 680 5261 686 5295
rect 504 5223 686 5261
rect 504 5189 646 5223
rect 680 5189 686 5223
rect 504 5151 686 5189
rect 504 5117 646 5151
rect 680 5117 686 5151
rect 504 5079 686 5117
rect 504 5045 646 5079
rect 680 5045 686 5079
rect 504 5007 686 5045
rect 504 4973 646 5007
rect 680 4973 686 5007
rect 504 4935 686 4973
rect 504 4901 646 4935
rect 680 4901 686 4935
rect 504 4863 686 4901
rect 504 4829 646 4863
rect 680 4829 686 4863
rect 504 4791 686 4829
rect 504 4757 646 4791
rect 680 4757 686 4791
rect 504 4719 686 4757
rect 504 4685 646 4719
rect 680 4685 686 4719
rect 504 4647 686 4685
rect 504 4613 646 4647
rect 680 4613 686 4647
rect 504 4575 686 4613
rect 504 4541 646 4575
rect 680 4541 686 4575
rect 504 4503 686 4541
rect 504 4469 646 4503
rect 680 4469 686 4503
rect 504 4431 686 4469
rect 504 4397 646 4431
rect 680 4397 686 4431
rect 504 4359 686 4397
rect 504 4325 646 4359
rect 680 4325 686 4359
rect 504 4287 686 4325
rect 504 4253 646 4287
rect 680 4253 686 4287
rect 504 4215 686 4253
rect 504 4181 646 4215
rect 680 4181 686 4215
rect 504 4143 686 4181
rect 504 4109 646 4143
rect 680 4109 686 4143
rect 504 4071 686 4109
rect 504 4037 646 4071
rect 680 4037 686 4071
rect 504 3999 686 4037
rect 504 3965 646 3999
rect 680 3965 686 3999
rect 504 3927 686 3965
rect 504 3893 646 3927
rect 680 3893 686 3927
rect 504 3855 686 3893
rect 504 3821 646 3855
rect 680 3821 686 3855
rect 504 3783 686 3821
rect 504 3749 646 3783
rect 680 3749 686 3783
rect 504 3711 686 3749
rect 504 3677 646 3711
rect 680 3677 686 3711
rect 504 3630 686 3677
rect 898 5583 1080 5630
rect 898 5549 904 5583
rect 938 5549 1080 5583
rect 898 5511 1080 5549
rect 898 5477 904 5511
rect 938 5477 1080 5511
rect 898 5439 1080 5477
rect 898 5405 904 5439
rect 938 5405 1080 5439
rect 898 5367 1080 5405
rect 898 5333 904 5367
rect 938 5333 1080 5367
rect 898 5295 1080 5333
rect 898 5261 904 5295
rect 938 5261 1080 5295
rect 898 5223 1080 5261
rect 898 5189 904 5223
rect 938 5189 1080 5223
rect 898 5151 1080 5189
rect 898 5117 904 5151
rect 938 5117 1080 5151
rect 898 5079 1080 5117
rect 898 5045 904 5079
rect 938 5045 1080 5079
rect 898 5007 1080 5045
rect 898 4973 904 5007
rect 938 4973 1080 5007
rect 898 4935 1080 4973
rect 898 4901 904 4935
rect 938 4901 1080 4935
rect 898 4863 1080 4901
rect 898 4829 904 4863
rect 938 4829 1080 4863
rect 898 4791 1080 4829
rect 898 4757 904 4791
rect 938 4757 1080 4791
rect 898 4719 1080 4757
rect 898 4685 904 4719
rect 938 4685 1080 4719
rect 898 4647 1080 4685
rect 898 4613 904 4647
rect 938 4613 1080 4647
rect 898 4575 1080 4613
rect 898 4541 904 4575
rect 938 4541 1080 4575
rect 898 4503 1080 4541
rect 898 4469 904 4503
rect 938 4469 1080 4503
rect 898 4431 1080 4469
rect 898 4397 904 4431
rect 938 4397 1080 4431
rect 898 4359 1080 4397
rect 898 4325 904 4359
rect 938 4325 1080 4359
rect 898 4287 1080 4325
rect 898 4253 904 4287
rect 938 4253 1080 4287
rect 898 4215 1080 4253
rect 898 4181 904 4215
rect 938 4181 1080 4215
rect 898 4143 1080 4181
rect 898 4109 904 4143
rect 938 4109 1080 4143
rect 898 4071 1080 4109
rect 898 4037 904 4071
rect 938 4037 1080 4071
rect 898 3999 1080 4037
rect 898 3965 904 3999
rect 938 3965 1080 3999
rect 898 3927 1080 3965
rect 898 3893 904 3927
rect 938 3893 1080 3927
rect 898 3855 1080 3893
rect 898 3821 904 3855
rect 938 3821 1080 3855
rect 898 3783 1080 3821
rect 898 3749 904 3783
rect 938 3749 1080 3783
rect 898 3711 1080 3749
rect 898 3677 904 3711
rect 938 3677 1080 3711
rect 898 3630 1080 3677
rect 1204 5583 1386 5630
rect 1204 5549 1346 5583
rect 1380 5549 1386 5583
rect 1204 5511 1386 5549
rect 1204 5477 1346 5511
rect 1380 5477 1386 5511
rect 1204 5439 1386 5477
rect 1204 5405 1346 5439
rect 1380 5405 1386 5439
rect 1204 5367 1386 5405
rect 1204 5333 1346 5367
rect 1380 5333 1386 5367
rect 1204 5295 1386 5333
rect 1204 5261 1346 5295
rect 1380 5261 1386 5295
rect 1204 5223 1386 5261
rect 1204 5189 1346 5223
rect 1380 5189 1386 5223
rect 1204 5151 1386 5189
rect 1204 5117 1346 5151
rect 1380 5117 1386 5151
rect 1204 5079 1386 5117
rect 1204 5045 1346 5079
rect 1380 5045 1386 5079
rect 1204 5007 1386 5045
rect 1204 4973 1346 5007
rect 1380 4973 1386 5007
rect 1204 4935 1386 4973
rect 1204 4901 1346 4935
rect 1380 4901 1386 4935
rect 1204 4863 1386 4901
rect 1204 4829 1346 4863
rect 1380 4829 1386 4863
rect 1204 4791 1386 4829
rect 1204 4757 1346 4791
rect 1380 4757 1386 4791
rect 1204 4719 1386 4757
rect 1204 4685 1346 4719
rect 1380 4685 1386 4719
rect 1204 4647 1386 4685
rect 1204 4613 1346 4647
rect 1380 4613 1386 4647
rect 1204 4575 1386 4613
rect 1204 4541 1346 4575
rect 1380 4541 1386 4575
rect 1204 4503 1386 4541
rect 1204 4469 1346 4503
rect 1380 4469 1386 4503
rect 1204 4431 1386 4469
rect 1204 4397 1346 4431
rect 1380 4397 1386 4431
rect 1204 4359 1386 4397
rect 1204 4325 1346 4359
rect 1380 4325 1386 4359
rect 1204 4287 1386 4325
rect 1204 4253 1346 4287
rect 1380 4253 1386 4287
rect 1204 4215 1386 4253
rect 1204 4181 1346 4215
rect 1380 4181 1386 4215
rect 1204 4143 1386 4181
rect 1204 4109 1346 4143
rect 1380 4109 1386 4143
rect 1204 4071 1386 4109
rect 1204 4037 1346 4071
rect 1380 4037 1386 4071
rect 1204 3999 1386 4037
rect 1204 3965 1346 3999
rect 1380 3965 1386 3999
rect 1204 3927 1386 3965
rect 1204 3893 1346 3927
rect 1380 3893 1386 3927
rect 1204 3855 1386 3893
rect 1204 3821 1346 3855
rect 1380 3821 1386 3855
rect 1204 3783 1386 3821
rect 1204 3749 1346 3783
rect 1380 3749 1386 3783
rect 1204 3711 1386 3749
rect 1204 3677 1346 3711
rect 1380 3677 1386 3711
rect 1204 3630 1386 3677
rect 1598 5583 1780 5630
rect 1598 5549 1604 5583
rect 1638 5549 1780 5583
rect 1598 5511 1780 5549
rect 1598 5477 1604 5511
rect 1638 5477 1780 5511
rect 1598 5439 1780 5477
rect 1598 5405 1604 5439
rect 1638 5405 1780 5439
rect 1598 5367 1780 5405
rect 1598 5333 1604 5367
rect 1638 5333 1780 5367
rect 1598 5295 1780 5333
rect 1598 5261 1604 5295
rect 1638 5261 1780 5295
rect 1598 5223 1780 5261
rect 1598 5189 1604 5223
rect 1638 5189 1780 5223
rect 1598 5151 1780 5189
rect 1598 5117 1604 5151
rect 1638 5117 1780 5151
rect 1598 5079 1780 5117
rect 1598 5045 1604 5079
rect 1638 5045 1780 5079
rect 1598 5007 1780 5045
rect 1598 4973 1604 5007
rect 1638 4973 1780 5007
rect 1598 4935 1780 4973
rect 1598 4901 1604 4935
rect 1638 4901 1780 4935
rect 1598 4863 1780 4901
rect 1598 4829 1604 4863
rect 1638 4829 1780 4863
rect 1598 4791 1780 4829
rect 1598 4757 1604 4791
rect 1638 4757 1780 4791
rect 1598 4719 1780 4757
rect 1598 4685 1604 4719
rect 1638 4685 1780 4719
rect 1598 4647 1780 4685
rect 1598 4613 1604 4647
rect 1638 4613 1780 4647
rect 1598 4575 1780 4613
rect 1598 4541 1604 4575
rect 1638 4541 1780 4575
rect 1598 4503 1780 4541
rect 1598 4469 1604 4503
rect 1638 4469 1780 4503
rect 1598 4431 1780 4469
rect 1598 4397 1604 4431
rect 1638 4397 1780 4431
rect 1598 4359 1780 4397
rect 1598 4325 1604 4359
rect 1638 4325 1780 4359
rect 1598 4287 1780 4325
rect 1598 4253 1604 4287
rect 1638 4253 1780 4287
rect 1598 4215 1780 4253
rect 1598 4181 1604 4215
rect 1638 4181 1780 4215
rect 1598 4143 1780 4181
rect 1598 4109 1604 4143
rect 1638 4109 1780 4143
rect 1598 4071 1780 4109
rect 1598 4037 1604 4071
rect 1638 4037 1780 4071
rect 1598 3999 1780 4037
rect 1598 3965 1604 3999
rect 1638 3965 1780 3999
rect 1598 3927 1780 3965
rect 1598 3893 1604 3927
rect 1638 3893 1780 3927
rect 1598 3855 1780 3893
rect 1598 3821 1604 3855
rect 1638 3821 1780 3855
rect 1598 3783 1780 3821
rect 1598 3749 1604 3783
rect 1638 3749 1780 3783
rect 1598 3711 1780 3749
rect 1598 3677 1604 3711
rect 1638 3677 1780 3711
rect 1598 3630 1780 3677
rect 1904 5583 2086 5630
rect 1904 5549 2046 5583
rect 2080 5549 2086 5583
rect 1904 5511 2086 5549
rect 1904 5477 2046 5511
rect 2080 5477 2086 5511
rect 1904 5439 2086 5477
rect 1904 5405 2046 5439
rect 2080 5405 2086 5439
rect 1904 5367 2086 5405
rect 1904 5333 2046 5367
rect 2080 5333 2086 5367
rect 1904 5295 2086 5333
rect 1904 5261 2046 5295
rect 2080 5261 2086 5295
rect 1904 5223 2086 5261
rect 1904 5189 2046 5223
rect 2080 5189 2086 5223
rect 1904 5151 2086 5189
rect 1904 5117 2046 5151
rect 2080 5117 2086 5151
rect 1904 5079 2086 5117
rect 1904 5045 2046 5079
rect 2080 5045 2086 5079
rect 1904 5007 2086 5045
rect 1904 4973 2046 5007
rect 2080 4973 2086 5007
rect 1904 4935 2086 4973
rect 1904 4901 2046 4935
rect 2080 4901 2086 4935
rect 1904 4863 2086 4901
rect 1904 4829 2046 4863
rect 2080 4829 2086 4863
rect 1904 4791 2086 4829
rect 1904 4757 2046 4791
rect 2080 4757 2086 4791
rect 1904 4719 2086 4757
rect 1904 4685 2046 4719
rect 2080 4685 2086 4719
rect 1904 4647 2086 4685
rect 1904 4613 2046 4647
rect 2080 4613 2086 4647
rect 1904 4575 2086 4613
rect 1904 4541 2046 4575
rect 2080 4541 2086 4575
rect 1904 4503 2086 4541
rect 1904 4469 2046 4503
rect 2080 4469 2086 4503
rect 1904 4431 2086 4469
rect 1904 4397 2046 4431
rect 2080 4397 2086 4431
rect 1904 4359 2086 4397
rect 1904 4325 2046 4359
rect 2080 4325 2086 4359
rect 1904 4287 2086 4325
rect 1904 4253 2046 4287
rect 2080 4253 2086 4287
rect 1904 4215 2086 4253
rect 1904 4181 2046 4215
rect 2080 4181 2086 4215
rect 1904 4143 2086 4181
rect 1904 4109 2046 4143
rect 2080 4109 2086 4143
rect 1904 4071 2086 4109
rect 1904 4037 2046 4071
rect 2080 4037 2086 4071
rect 1904 3999 2086 4037
rect 1904 3965 2046 3999
rect 2080 3965 2086 3999
rect 1904 3927 2086 3965
rect 1904 3893 2046 3927
rect 2080 3893 2086 3927
rect 1904 3855 2086 3893
rect 1904 3821 2046 3855
rect 2080 3821 2086 3855
rect 1904 3783 2086 3821
rect 1904 3749 2046 3783
rect 2080 3749 2086 3783
rect 1904 3711 2086 3749
rect 1904 3677 2046 3711
rect 2080 3677 2086 3711
rect 1904 3630 2086 3677
rect 2298 5583 2480 5630
rect 2298 5549 2304 5583
rect 2338 5549 2480 5583
rect 2298 5511 2480 5549
rect 2298 5477 2304 5511
rect 2338 5477 2480 5511
rect 2298 5439 2480 5477
rect 2298 5405 2304 5439
rect 2338 5405 2480 5439
rect 2298 5367 2480 5405
rect 2298 5333 2304 5367
rect 2338 5333 2480 5367
rect 2298 5295 2480 5333
rect 2298 5261 2304 5295
rect 2338 5261 2480 5295
rect 2298 5223 2480 5261
rect 2298 5189 2304 5223
rect 2338 5189 2480 5223
rect 2298 5151 2480 5189
rect 2298 5117 2304 5151
rect 2338 5117 2480 5151
rect 2298 5079 2480 5117
rect 2298 5045 2304 5079
rect 2338 5045 2480 5079
rect 2298 5007 2480 5045
rect 2298 4973 2304 5007
rect 2338 4973 2480 5007
rect 2298 4935 2480 4973
rect 2298 4901 2304 4935
rect 2338 4901 2480 4935
rect 2298 4863 2480 4901
rect 2298 4829 2304 4863
rect 2338 4829 2480 4863
rect 2298 4791 2480 4829
rect 2298 4757 2304 4791
rect 2338 4757 2480 4791
rect 2298 4719 2480 4757
rect 2298 4685 2304 4719
rect 2338 4685 2480 4719
rect 2298 4647 2480 4685
rect 2298 4613 2304 4647
rect 2338 4613 2480 4647
rect 2298 4575 2480 4613
rect 2298 4541 2304 4575
rect 2338 4541 2480 4575
rect 2298 4503 2480 4541
rect 2298 4469 2304 4503
rect 2338 4469 2480 4503
rect 2298 4431 2480 4469
rect 2298 4397 2304 4431
rect 2338 4397 2480 4431
rect 2298 4359 2480 4397
rect 2298 4325 2304 4359
rect 2338 4325 2480 4359
rect 2298 4287 2480 4325
rect 2298 4253 2304 4287
rect 2338 4253 2480 4287
rect 2298 4215 2480 4253
rect 2298 4181 2304 4215
rect 2338 4181 2480 4215
rect 2298 4143 2480 4181
rect 2298 4109 2304 4143
rect 2338 4109 2480 4143
rect 2298 4071 2480 4109
rect 2298 4037 2304 4071
rect 2338 4037 2480 4071
rect 2298 3999 2480 4037
rect 2298 3965 2304 3999
rect 2338 3965 2480 3999
rect 2298 3927 2480 3965
rect 2298 3893 2304 3927
rect 2338 3893 2480 3927
rect 2298 3855 2480 3893
rect 2298 3821 2304 3855
rect 2338 3821 2480 3855
rect 2298 3783 2480 3821
rect 2298 3749 2304 3783
rect 2338 3749 2480 3783
rect 2298 3711 2480 3749
rect 2298 3677 2304 3711
rect 2338 3677 2480 3711
rect 2298 3630 2480 3677
rect 3604 5583 3786 5630
rect 3604 5549 3746 5583
rect 3780 5549 3786 5583
rect 3604 5511 3786 5549
rect 3604 5477 3746 5511
rect 3780 5477 3786 5511
rect 3604 5439 3786 5477
rect 3604 5405 3746 5439
rect 3780 5405 3786 5439
rect 3604 5367 3786 5405
rect 3604 5333 3746 5367
rect 3780 5333 3786 5367
rect 3604 5295 3786 5333
rect 3604 5261 3746 5295
rect 3780 5261 3786 5295
rect 3604 5223 3786 5261
rect 3604 5189 3746 5223
rect 3780 5189 3786 5223
rect 3604 5151 3786 5189
rect 3604 5117 3746 5151
rect 3780 5117 3786 5151
rect 3604 5079 3786 5117
rect 3604 5045 3746 5079
rect 3780 5045 3786 5079
rect 3604 5007 3786 5045
rect 3604 4973 3746 5007
rect 3780 4973 3786 5007
rect 3604 4935 3786 4973
rect 3604 4901 3746 4935
rect 3780 4901 3786 4935
rect 3604 4863 3786 4901
rect 3604 4829 3746 4863
rect 3780 4829 3786 4863
rect 3604 4791 3786 4829
rect 3604 4757 3746 4791
rect 3780 4757 3786 4791
rect 3604 4719 3786 4757
rect 3604 4685 3746 4719
rect 3780 4685 3786 4719
rect 3604 4647 3786 4685
rect 3604 4613 3746 4647
rect 3780 4613 3786 4647
rect 3604 4575 3786 4613
rect 3604 4541 3746 4575
rect 3780 4541 3786 4575
rect 3604 4503 3786 4541
rect 3604 4469 3746 4503
rect 3780 4469 3786 4503
rect 3604 4431 3786 4469
rect 3604 4397 3746 4431
rect 3780 4397 3786 4431
rect 3604 4359 3786 4397
rect 3604 4325 3746 4359
rect 3780 4325 3786 4359
rect 3604 4287 3786 4325
rect 3604 4253 3746 4287
rect 3780 4253 3786 4287
rect 3604 4215 3786 4253
rect 3604 4181 3746 4215
rect 3780 4181 3786 4215
rect 3604 4143 3786 4181
rect 3604 4109 3746 4143
rect 3780 4109 3786 4143
rect 3604 4071 3786 4109
rect 3604 4037 3746 4071
rect 3780 4037 3786 4071
rect 3604 3999 3786 4037
rect 3604 3965 3746 3999
rect 3780 3965 3786 3999
rect 3604 3927 3786 3965
rect 3604 3893 3746 3927
rect 3780 3893 3786 3927
rect 3604 3855 3786 3893
rect 3604 3821 3746 3855
rect 3780 3821 3786 3855
rect 3604 3783 3786 3821
rect 3604 3749 3746 3783
rect 3780 3749 3786 3783
rect 3604 3711 3786 3749
rect 3604 3677 3746 3711
rect 3780 3677 3786 3711
rect 3604 3630 3786 3677
rect 3998 5583 4180 5630
rect 3998 5549 4004 5583
rect 4038 5549 4180 5583
rect 3998 5511 4180 5549
rect 3998 5477 4004 5511
rect 4038 5477 4180 5511
rect 3998 5439 4180 5477
rect 3998 5405 4004 5439
rect 4038 5405 4180 5439
rect 3998 5367 4180 5405
rect 3998 5333 4004 5367
rect 4038 5333 4180 5367
rect 3998 5295 4180 5333
rect 3998 5261 4004 5295
rect 4038 5261 4180 5295
rect 3998 5223 4180 5261
rect 3998 5189 4004 5223
rect 4038 5189 4180 5223
rect 3998 5151 4180 5189
rect 3998 5117 4004 5151
rect 4038 5117 4180 5151
rect 3998 5079 4180 5117
rect 3998 5045 4004 5079
rect 4038 5045 4180 5079
rect 3998 5007 4180 5045
rect 3998 4973 4004 5007
rect 4038 4973 4180 5007
rect 3998 4935 4180 4973
rect 3998 4901 4004 4935
rect 4038 4901 4180 4935
rect 3998 4863 4180 4901
rect 3998 4829 4004 4863
rect 4038 4829 4180 4863
rect 3998 4791 4180 4829
rect 3998 4757 4004 4791
rect 4038 4757 4180 4791
rect 3998 4719 4180 4757
rect 3998 4685 4004 4719
rect 4038 4685 4180 4719
rect 3998 4647 4180 4685
rect 3998 4613 4004 4647
rect 4038 4613 4180 4647
rect 3998 4575 4180 4613
rect 3998 4541 4004 4575
rect 4038 4541 4180 4575
rect 3998 4503 4180 4541
rect 3998 4469 4004 4503
rect 4038 4469 4180 4503
rect 3998 4431 4180 4469
rect 3998 4397 4004 4431
rect 4038 4397 4180 4431
rect 3998 4359 4180 4397
rect 3998 4325 4004 4359
rect 4038 4325 4180 4359
rect 3998 4287 4180 4325
rect 3998 4253 4004 4287
rect 4038 4253 4180 4287
rect 3998 4215 4180 4253
rect 3998 4181 4004 4215
rect 4038 4181 4180 4215
rect 3998 4143 4180 4181
rect 3998 4109 4004 4143
rect 4038 4109 4180 4143
rect 3998 4071 4180 4109
rect 3998 4037 4004 4071
rect 4038 4037 4180 4071
rect 3998 3999 4180 4037
rect 3998 3965 4004 3999
rect 4038 3965 4180 3999
rect 3998 3927 4180 3965
rect 3998 3893 4004 3927
rect 4038 3893 4180 3927
rect 3998 3855 4180 3893
rect 3998 3821 4004 3855
rect 4038 3821 4180 3855
rect 3998 3783 4180 3821
rect 3998 3749 4004 3783
rect 4038 3749 4180 3783
rect 3998 3711 4180 3749
rect 3998 3677 4004 3711
rect 4038 3677 4180 3711
rect 3998 3630 4180 3677
rect 4304 5583 4486 5630
rect 4304 5549 4446 5583
rect 4480 5549 4486 5583
rect 4304 5511 4486 5549
rect 4304 5477 4446 5511
rect 4480 5477 4486 5511
rect 4304 5439 4486 5477
rect 4304 5405 4446 5439
rect 4480 5405 4486 5439
rect 4304 5367 4486 5405
rect 4304 5333 4446 5367
rect 4480 5333 4486 5367
rect 4304 5295 4486 5333
rect 4304 5261 4446 5295
rect 4480 5261 4486 5295
rect 4304 5223 4486 5261
rect 4304 5189 4446 5223
rect 4480 5189 4486 5223
rect 4304 5151 4486 5189
rect 4304 5117 4446 5151
rect 4480 5117 4486 5151
rect 4304 5079 4486 5117
rect 4304 5045 4446 5079
rect 4480 5045 4486 5079
rect 4304 5007 4486 5045
rect 4304 4973 4446 5007
rect 4480 4973 4486 5007
rect 4304 4935 4486 4973
rect 4304 4901 4446 4935
rect 4480 4901 4486 4935
rect 4304 4863 4486 4901
rect 4304 4829 4446 4863
rect 4480 4829 4486 4863
rect 4304 4791 4486 4829
rect 4304 4757 4446 4791
rect 4480 4757 4486 4791
rect 4304 4719 4486 4757
rect 4304 4685 4446 4719
rect 4480 4685 4486 4719
rect 4304 4647 4486 4685
rect 4304 4613 4446 4647
rect 4480 4613 4486 4647
rect 4304 4575 4486 4613
rect 4304 4541 4446 4575
rect 4480 4541 4486 4575
rect 4304 4503 4486 4541
rect 4304 4469 4446 4503
rect 4480 4469 4486 4503
rect 4304 4431 4486 4469
rect 4304 4397 4446 4431
rect 4480 4397 4486 4431
rect 4304 4359 4486 4397
rect 4304 4325 4446 4359
rect 4480 4325 4486 4359
rect 4304 4287 4486 4325
rect 4304 4253 4446 4287
rect 4480 4253 4486 4287
rect 4304 4215 4486 4253
rect 4304 4181 4446 4215
rect 4480 4181 4486 4215
rect 4304 4143 4486 4181
rect 4304 4109 4446 4143
rect 4480 4109 4486 4143
rect 4304 4071 4486 4109
rect 4304 4037 4446 4071
rect 4480 4037 4486 4071
rect 4304 3999 4486 4037
rect 4304 3965 4446 3999
rect 4480 3965 4486 3999
rect 4304 3927 4486 3965
rect 4304 3893 4446 3927
rect 4480 3893 4486 3927
rect 4304 3855 4486 3893
rect 4304 3821 4446 3855
rect 4480 3821 4486 3855
rect 4304 3783 4486 3821
rect 4304 3749 4446 3783
rect 4480 3749 4486 3783
rect 4304 3711 4486 3749
rect 4304 3677 4446 3711
rect 4480 3677 4486 3711
rect 4304 3630 4486 3677
rect 4698 5583 4880 5630
rect 4698 5549 4704 5583
rect 4738 5549 4880 5583
rect 4698 5511 4880 5549
rect 4698 5477 4704 5511
rect 4738 5477 4880 5511
rect 4698 5439 4880 5477
rect 4698 5405 4704 5439
rect 4738 5405 4880 5439
rect 4698 5367 4880 5405
rect 4698 5333 4704 5367
rect 4738 5333 4880 5367
rect 4698 5295 4880 5333
rect 4698 5261 4704 5295
rect 4738 5261 4880 5295
rect 4698 5223 4880 5261
rect 4698 5189 4704 5223
rect 4738 5189 4880 5223
rect 4698 5151 4880 5189
rect 4698 5117 4704 5151
rect 4738 5117 4880 5151
rect 4698 5079 4880 5117
rect 4698 5045 4704 5079
rect 4738 5045 4880 5079
rect 4698 5007 4880 5045
rect 4698 4973 4704 5007
rect 4738 4973 4880 5007
rect 4698 4935 4880 4973
rect 4698 4901 4704 4935
rect 4738 4901 4880 4935
rect 4698 4863 4880 4901
rect 4698 4829 4704 4863
rect 4738 4829 4880 4863
rect 4698 4791 4880 4829
rect 4698 4757 4704 4791
rect 4738 4757 4880 4791
rect 4698 4719 4880 4757
rect 4698 4685 4704 4719
rect 4738 4685 4880 4719
rect 4698 4647 4880 4685
rect 4698 4613 4704 4647
rect 4738 4613 4880 4647
rect 4698 4575 4880 4613
rect 4698 4541 4704 4575
rect 4738 4541 4880 4575
rect 4698 4503 4880 4541
rect 4698 4469 4704 4503
rect 4738 4469 4880 4503
rect 4698 4431 4880 4469
rect 4698 4397 4704 4431
rect 4738 4397 4880 4431
rect 4698 4359 4880 4397
rect 4698 4325 4704 4359
rect 4738 4325 4880 4359
rect 4698 4287 4880 4325
rect 4698 4253 4704 4287
rect 4738 4253 4880 4287
rect 4698 4215 4880 4253
rect 4698 4181 4704 4215
rect 4738 4181 4880 4215
rect 4698 4143 4880 4181
rect 4698 4109 4704 4143
rect 4738 4109 4880 4143
rect 4698 4071 4880 4109
rect 4698 4037 4704 4071
rect 4738 4037 4880 4071
rect 4698 3999 4880 4037
rect 4698 3965 4704 3999
rect 4738 3965 4880 3999
rect 4698 3927 4880 3965
rect 4698 3893 4704 3927
rect 4738 3893 4880 3927
rect 4698 3855 4880 3893
rect 4698 3821 4704 3855
rect 4738 3821 4880 3855
rect 4698 3783 4880 3821
rect 4698 3749 4704 3783
rect 4738 3749 4880 3783
rect 4698 3711 4880 3749
rect 4698 3677 4704 3711
rect 4738 3677 4880 3711
rect 4698 3630 4880 3677
rect 5004 5583 5186 5630
rect 5004 5549 5146 5583
rect 5180 5549 5186 5583
rect 5004 5511 5186 5549
rect 5004 5477 5146 5511
rect 5180 5477 5186 5511
rect 5004 5439 5186 5477
rect 5004 5405 5146 5439
rect 5180 5405 5186 5439
rect 5004 5367 5186 5405
rect 5004 5333 5146 5367
rect 5180 5333 5186 5367
rect 5004 5295 5186 5333
rect 5004 5261 5146 5295
rect 5180 5261 5186 5295
rect 5004 5223 5186 5261
rect 5004 5189 5146 5223
rect 5180 5189 5186 5223
rect 5004 5151 5186 5189
rect 5004 5117 5146 5151
rect 5180 5117 5186 5151
rect 5004 5079 5186 5117
rect 5004 5045 5146 5079
rect 5180 5045 5186 5079
rect 5004 5007 5186 5045
rect 5004 4973 5146 5007
rect 5180 4973 5186 5007
rect 5004 4935 5186 4973
rect 5004 4901 5146 4935
rect 5180 4901 5186 4935
rect 5004 4863 5186 4901
rect 5004 4829 5146 4863
rect 5180 4829 5186 4863
rect 5004 4791 5186 4829
rect 5004 4757 5146 4791
rect 5180 4757 5186 4791
rect 5004 4719 5186 4757
rect 5004 4685 5146 4719
rect 5180 4685 5186 4719
rect 5004 4647 5186 4685
rect 5004 4613 5146 4647
rect 5180 4613 5186 4647
rect 5004 4575 5186 4613
rect 5004 4541 5146 4575
rect 5180 4541 5186 4575
rect 5004 4503 5186 4541
rect 5004 4469 5146 4503
rect 5180 4469 5186 4503
rect 5004 4431 5186 4469
rect 5004 4397 5146 4431
rect 5180 4397 5186 4431
rect 5004 4359 5186 4397
rect 5004 4325 5146 4359
rect 5180 4325 5186 4359
rect 5004 4287 5186 4325
rect 5004 4253 5146 4287
rect 5180 4253 5186 4287
rect 5004 4215 5186 4253
rect 5004 4181 5146 4215
rect 5180 4181 5186 4215
rect 5004 4143 5186 4181
rect 5004 4109 5146 4143
rect 5180 4109 5186 4143
rect 5004 4071 5186 4109
rect 5004 4037 5146 4071
rect 5180 4037 5186 4071
rect 5004 3999 5186 4037
rect 5004 3965 5146 3999
rect 5180 3965 5186 3999
rect 5004 3927 5186 3965
rect 5004 3893 5146 3927
rect 5180 3893 5186 3927
rect 5004 3855 5186 3893
rect 5004 3821 5146 3855
rect 5180 3821 5186 3855
rect 5004 3783 5186 3821
rect 5004 3749 5146 3783
rect 5180 3749 5186 3783
rect 5004 3711 5186 3749
rect 5004 3677 5146 3711
rect 5180 3677 5186 3711
rect 5004 3630 5186 3677
rect 5398 5583 5580 5630
rect 5398 5549 5404 5583
rect 5438 5549 5580 5583
rect 5398 5511 5580 5549
rect 5398 5477 5404 5511
rect 5438 5477 5580 5511
rect 5398 5439 5580 5477
rect 5398 5405 5404 5439
rect 5438 5405 5580 5439
rect 5398 5367 5580 5405
rect 5398 5333 5404 5367
rect 5438 5333 5580 5367
rect 5398 5295 5580 5333
rect 5398 5261 5404 5295
rect 5438 5261 5580 5295
rect 5398 5223 5580 5261
rect 5398 5189 5404 5223
rect 5438 5189 5580 5223
rect 5398 5151 5580 5189
rect 5398 5117 5404 5151
rect 5438 5117 5580 5151
rect 5398 5079 5580 5117
rect 5398 5045 5404 5079
rect 5438 5045 5580 5079
rect 5398 5007 5580 5045
rect 5398 4973 5404 5007
rect 5438 4973 5580 5007
rect 5398 4935 5580 4973
rect 5398 4901 5404 4935
rect 5438 4901 5580 4935
rect 5398 4863 5580 4901
rect 5398 4829 5404 4863
rect 5438 4829 5580 4863
rect 5398 4791 5580 4829
rect 5398 4757 5404 4791
rect 5438 4757 5580 4791
rect 5398 4719 5580 4757
rect 5398 4685 5404 4719
rect 5438 4685 5580 4719
rect 5398 4647 5580 4685
rect 5398 4613 5404 4647
rect 5438 4613 5580 4647
rect 5398 4575 5580 4613
rect 5398 4541 5404 4575
rect 5438 4541 5580 4575
rect 5398 4503 5580 4541
rect 5398 4469 5404 4503
rect 5438 4469 5580 4503
rect 5398 4431 5580 4469
rect 5398 4397 5404 4431
rect 5438 4397 5580 4431
rect 5398 4359 5580 4397
rect 5398 4325 5404 4359
rect 5438 4325 5580 4359
rect 5398 4287 5580 4325
rect 5398 4253 5404 4287
rect 5438 4253 5580 4287
rect 5398 4215 5580 4253
rect 5398 4181 5404 4215
rect 5438 4181 5580 4215
rect 5398 4143 5580 4181
rect 5398 4109 5404 4143
rect 5438 4109 5580 4143
rect 5398 4071 5580 4109
rect 5398 4037 5404 4071
rect 5438 4037 5580 4071
rect 5398 3999 5580 4037
rect 5398 3965 5404 3999
rect 5438 3965 5580 3999
rect 5398 3927 5580 3965
rect 5398 3893 5404 3927
rect 5438 3893 5580 3927
rect 5398 3855 5580 3893
rect 5398 3821 5404 3855
rect 5438 3821 5580 3855
rect 5398 3783 5580 3821
rect 5398 3749 5404 3783
rect 5438 3749 5580 3783
rect 5398 3711 5580 3749
rect 5398 3677 5404 3711
rect 5438 3677 5580 3711
rect 5398 3630 5580 3677
rect 5704 5583 5886 5630
rect 5704 5549 5846 5583
rect 5880 5549 5886 5583
rect 5704 5511 5886 5549
rect 5704 5477 5846 5511
rect 5880 5477 5886 5511
rect 5704 5439 5886 5477
rect 5704 5405 5846 5439
rect 5880 5405 5886 5439
rect 5704 5367 5886 5405
rect 5704 5333 5846 5367
rect 5880 5333 5886 5367
rect 5704 5295 5886 5333
rect 5704 5261 5846 5295
rect 5880 5261 5886 5295
rect 5704 5223 5886 5261
rect 5704 5189 5846 5223
rect 5880 5189 5886 5223
rect 5704 5151 5886 5189
rect 5704 5117 5846 5151
rect 5880 5117 5886 5151
rect 5704 5079 5886 5117
rect 5704 5045 5846 5079
rect 5880 5045 5886 5079
rect 5704 5007 5886 5045
rect 5704 4973 5846 5007
rect 5880 4973 5886 5007
rect 5704 4935 5886 4973
rect 5704 4901 5846 4935
rect 5880 4901 5886 4935
rect 5704 4863 5886 4901
rect 5704 4829 5846 4863
rect 5880 4829 5886 4863
rect 5704 4791 5886 4829
rect 5704 4757 5846 4791
rect 5880 4757 5886 4791
rect 5704 4719 5886 4757
rect 5704 4685 5846 4719
rect 5880 4685 5886 4719
rect 5704 4647 5886 4685
rect 5704 4613 5846 4647
rect 5880 4613 5886 4647
rect 5704 4575 5886 4613
rect 5704 4541 5846 4575
rect 5880 4541 5886 4575
rect 5704 4503 5886 4541
rect 5704 4469 5846 4503
rect 5880 4469 5886 4503
rect 5704 4431 5886 4469
rect 5704 4397 5846 4431
rect 5880 4397 5886 4431
rect 5704 4359 5886 4397
rect 5704 4325 5846 4359
rect 5880 4325 5886 4359
rect 5704 4287 5886 4325
rect 5704 4253 5846 4287
rect 5880 4253 5886 4287
rect 5704 4215 5886 4253
rect 5704 4181 5846 4215
rect 5880 4181 5886 4215
rect 5704 4143 5886 4181
rect 5704 4109 5846 4143
rect 5880 4109 5886 4143
rect 5704 4071 5886 4109
rect 5704 4037 5846 4071
rect 5880 4037 5886 4071
rect 5704 3999 5886 4037
rect 5704 3965 5846 3999
rect 5880 3965 5886 3999
rect 5704 3927 5886 3965
rect 5704 3893 5846 3927
rect 5880 3893 5886 3927
rect 5704 3855 5886 3893
rect 5704 3821 5846 3855
rect 5880 3821 5886 3855
rect 5704 3783 5886 3821
rect 5704 3749 5846 3783
rect 5880 3749 5886 3783
rect 5704 3711 5886 3749
rect 5704 3677 5846 3711
rect 5880 3677 5886 3711
rect 5704 3630 5886 3677
rect 6098 5583 6280 5630
rect 6098 5549 6104 5583
rect 6138 5549 6280 5583
rect 6098 5511 6280 5549
rect 6098 5477 6104 5511
rect 6138 5477 6280 5511
rect 6098 5439 6280 5477
rect 6098 5405 6104 5439
rect 6138 5405 6280 5439
rect 6098 5367 6280 5405
rect 6098 5333 6104 5367
rect 6138 5333 6280 5367
rect 6098 5295 6280 5333
rect 6098 5261 6104 5295
rect 6138 5261 6280 5295
rect 6098 5223 6280 5261
rect 6098 5189 6104 5223
rect 6138 5189 6280 5223
rect 6098 5151 6280 5189
rect 6098 5117 6104 5151
rect 6138 5117 6280 5151
rect 6098 5079 6280 5117
rect 6098 5045 6104 5079
rect 6138 5045 6280 5079
rect 6098 5007 6280 5045
rect 6098 4973 6104 5007
rect 6138 4973 6280 5007
rect 6098 4935 6280 4973
rect 6098 4901 6104 4935
rect 6138 4901 6280 4935
rect 6098 4863 6280 4901
rect 6098 4829 6104 4863
rect 6138 4829 6280 4863
rect 6098 4791 6280 4829
rect 6098 4757 6104 4791
rect 6138 4757 6280 4791
rect 6098 4719 6280 4757
rect 6098 4685 6104 4719
rect 6138 4685 6280 4719
rect 6098 4647 6280 4685
rect 6098 4613 6104 4647
rect 6138 4613 6280 4647
rect 6098 4575 6280 4613
rect 6098 4541 6104 4575
rect 6138 4541 6280 4575
rect 6098 4503 6280 4541
rect 6098 4469 6104 4503
rect 6138 4469 6280 4503
rect 6098 4431 6280 4469
rect 6098 4397 6104 4431
rect 6138 4397 6280 4431
rect 6098 4359 6280 4397
rect 6098 4325 6104 4359
rect 6138 4325 6280 4359
rect 6098 4287 6280 4325
rect 6098 4253 6104 4287
rect 6138 4253 6280 4287
rect 6098 4215 6280 4253
rect 6098 4181 6104 4215
rect 6138 4181 6280 4215
rect 6098 4143 6280 4181
rect 6098 4109 6104 4143
rect 6138 4109 6280 4143
rect 6098 4071 6280 4109
rect 6098 4037 6104 4071
rect 6138 4037 6280 4071
rect 6098 3999 6280 4037
rect 6098 3965 6104 3999
rect 6138 3965 6280 3999
rect 6098 3927 6280 3965
rect 6098 3893 6104 3927
rect 6138 3893 6280 3927
rect 6098 3855 6280 3893
rect 6098 3821 6104 3855
rect 6138 3821 6280 3855
rect 6098 3783 6280 3821
rect 6098 3749 6104 3783
rect 6138 3749 6280 3783
rect 6098 3711 6280 3749
rect 6098 3677 6104 3711
rect 6138 3677 6280 3711
rect 6098 3630 6280 3677
rect 6404 5583 6586 5630
rect 6404 5549 6546 5583
rect 6580 5549 6586 5583
rect 6404 5511 6586 5549
rect 6404 5477 6546 5511
rect 6580 5477 6586 5511
rect 6404 5439 6586 5477
rect 6404 5405 6546 5439
rect 6580 5405 6586 5439
rect 6404 5367 6586 5405
rect 6404 5333 6546 5367
rect 6580 5333 6586 5367
rect 6404 5295 6586 5333
rect 6404 5261 6546 5295
rect 6580 5261 6586 5295
rect 6404 5223 6586 5261
rect 6404 5189 6546 5223
rect 6580 5189 6586 5223
rect 6404 5151 6586 5189
rect 6404 5117 6546 5151
rect 6580 5117 6586 5151
rect 6404 5079 6586 5117
rect 6404 5045 6546 5079
rect 6580 5045 6586 5079
rect 6404 5007 6586 5045
rect 6404 4973 6546 5007
rect 6580 4973 6586 5007
rect 6404 4935 6586 4973
rect 6404 4901 6546 4935
rect 6580 4901 6586 4935
rect 6404 4863 6586 4901
rect 6404 4829 6546 4863
rect 6580 4829 6586 4863
rect 6404 4791 6586 4829
rect 6404 4757 6546 4791
rect 6580 4757 6586 4791
rect 6404 4719 6586 4757
rect 6404 4685 6546 4719
rect 6580 4685 6586 4719
rect 6404 4647 6586 4685
rect 6404 4613 6546 4647
rect 6580 4613 6586 4647
rect 6404 4575 6586 4613
rect 6404 4541 6546 4575
rect 6580 4541 6586 4575
rect 6404 4503 6586 4541
rect 6404 4469 6546 4503
rect 6580 4469 6586 4503
rect 6404 4431 6586 4469
rect 6404 4397 6546 4431
rect 6580 4397 6586 4431
rect 6404 4359 6586 4397
rect 6404 4325 6546 4359
rect 6580 4325 6586 4359
rect 6404 4287 6586 4325
rect 6404 4253 6546 4287
rect 6580 4253 6586 4287
rect 6404 4215 6586 4253
rect 6404 4181 6546 4215
rect 6580 4181 6586 4215
rect 6404 4143 6586 4181
rect 6404 4109 6546 4143
rect 6580 4109 6586 4143
rect 6404 4071 6586 4109
rect 6404 4037 6546 4071
rect 6580 4037 6586 4071
rect 6404 3999 6586 4037
rect 6404 3965 6546 3999
rect 6580 3965 6586 3999
rect 6404 3927 6586 3965
rect 6404 3893 6546 3927
rect 6580 3893 6586 3927
rect 6404 3855 6586 3893
rect 6404 3821 6546 3855
rect 6580 3821 6586 3855
rect 6404 3783 6586 3821
rect 6404 3749 6546 3783
rect 6580 3749 6586 3783
rect 6404 3711 6586 3749
rect 6404 3677 6546 3711
rect 6580 3677 6586 3711
rect 6404 3630 6586 3677
rect 6798 5583 6980 5630
rect 6798 5549 6804 5583
rect 6838 5549 6980 5583
rect 6798 5511 6980 5549
rect 6798 5477 6804 5511
rect 6838 5477 6980 5511
rect 6798 5439 6980 5477
rect 6798 5405 6804 5439
rect 6838 5405 6980 5439
rect 6798 5367 6980 5405
rect 6798 5333 6804 5367
rect 6838 5333 6980 5367
rect 6798 5295 6980 5333
rect 6798 5261 6804 5295
rect 6838 5261 6980 5295
rect 6798 5223 6980 5261
rect 6798 5189 6804 5223
rect 6838 5189 6980 5223
rect 6798 5151 6980 5189
rect 6798 5117 6804 5151
rect 6838 5117 6980 5151
rect 6798 5079 6980 5117
rect 6798 5045 6804 5079
rect 6838 5045 6980 5079
rect 6798 5007 6980 5045
rect 6798 4973 6804 5007
rect 6838 4973 6980 5007
rect 6798 4935 6980 4973
rect 6798 4901 6804 4935
rect 6838 4901 6980 4935
rect 6798 4863 6980 4901
rect 6798 4829 6804 4863
rect 6838 4829 6980 4863
rect 6798 4791 6980 4829
rect 6798 4757 6804 4791
rect 6838 4757 6980 4791
rect 6798 4719 6980 4757
rect 6798 4685 6804 4719
rect 6838 4685 6980 4719
rect 6798 4647 6980 4685
rect 6798 4613 6804 4647
rect 6838 4613 6980 4647
rect 6798 4575 6980 4613
rect 6798 4541 6804 4575
rect 6838 4541 6980 4575
rect 6798 4503 6980 4541
rect 6798 4469 6804 4503
rect 6838 4469 6980 4503
rect 6798 4431 6980 4469
rect 6798 4397 6804 4431
rect 6838 4397 6980 4431
rect 6798 4359 6980 4397
rect 6798 4325 6804 4359
rect 6838 4325 6980 4359
rect 6798 4287 6980 4325
rect 6798 4253 6804 4287
rect 6838 4253 6980 4287
rect 6798 4215 6980 4253
rect 6798 4181 6804 4215
rect 6838 4181 6980 4215
rect 6798 4143 6980 4181
rect 6798 4109 6804 4143
rect 6838 4109 6980 4143
rect 6798 4071 6980 4109
rect 6798 4037 6804 4071
rect 6838 4037 6980 4071
rect 6798 3999 6980 4037
rect 6798 3965 6804 3999
rect 6838 3965 6980 3999
rect 6798 3927 6980 3965
rect 6798 3893 6804 3927
rect 6838 3893 6980 3927
rect 6798 3855 6980 3893
rect 6798 3821 6804 3855
rect 6838 3821 6980 3855
rect 6798 3783 6980 3821
rect 6798 3749 6804 3783
rect 6838 3749 6980 3783
rect 6798 3711 6980 3749
rect 6798 3677 6804 3711
rect 6838 3677 6980 3711
rect 6798 3630 6980 3677
rect 7104 5583 7286 5630
rect 7104 5549 7246 5583
rect 7280 5549 7286 5583
rect 7104 5511 7286 5549
rect 7104 5477 7246 5511
rect 7280 5477 7286 5511
rect 7104 5439 7286 5477
rect 7104 5405 7246 5439
rect 7280 5405 7286 5439
rect 7104 5367 7286 5405
rect 7104 5333 7246 5367
rect 7280 5333 7286 5367
rect 7104 5295 7286 5333
rect 7104 5261 7246 5295
rect 7280 5261 7286 5295
rect 7104 5223 7286 5261
rect 7104 5189 7246 5223
rect 7280 5189 7286 5223
rect 7104 5151 7286 5189
rect 7104 5117 7246 5151
rect 7280 5117 7286 5151
rect 7104 5079 7286 5117
rect 7104 5045 7246 5079
rect 7280 5045 7286 5079
rect 7104 5007 7286 5045
rect 7104 4973 7246 5007
rect 7280 4973 7286 5007
rect 7104 4935 7286 4973
rect 7104 4901 7246 4935
rect 7280 4901 7286 4935
rect 7104 4863 7286 4901
rect 7104 4829 7246 4863
rect 7280 4829 7286 4863
rect 7104 4791 7286 4829
rect 7104 4757 7246 4791
rect 7280 4757 7286 4791
rect 7104 4719 7286 4757
rect 7104 4685 7246 4719
rect 7280 4685 7286 4719
rect 7104 4647 7286 4685
rect 7104 4613 7246 4647
rect 7280 4613 7286 4647
rect 7104 4575 7286 4613
rect 7104 4541 7246 4575
rect 7280 4541 7286 4575
rect 7104 4503 7286 4541
rect 7104 4469 7246 4503
rect 7280 4469 7286 4503
rect 7104 4431 7286 4469
rect 7104 4397 7246 4431
rect 7280 4397 7286 4431
rect 7104 4359 7286 4397
rect 7104 4325 7246 4359
rect 7280 4325 7286 4359
rect 7104 4287 7286 4325
rect 7104 4253 7246 4287
rect 7280 4253 7286 4287
rect 7104 4215 7286 4253
rect 7104 4181 7246 4215
rect 7280 4181 7286 4215
rect 7104 4143 7286 4181
rect 7104 4109 7246 4143
rect 7280 4109 7286 4143
rect 7104 4071 7286 4109
rect 7104 4037 7246 4071
rect 7280 4037 7286 4071
rect 7104 3999 7286 4037
rect 7104 3965 7246 3999
rect 7280 3965 7286 3999
rect 7104 3927 7286 3965
rect 7104 3893 7246 3927
rect 7280 3893 7286 3927
rect 7104 3855 7286 3893
rect 7104 3821 7246 3855
rect 7280 3821 7286 3855
rect 7104 3783 7286 3821
rect 7104 3749 7246 3783
rect 7280 3749 7286 3783
rect 7104 3711 7286 3749
rect 7104 3677 7246 3711
rect 7280 3677 7286 3711
rect 7104 3630 7286 3677
rect 7498 5583 7680 5630
rect 7498 5549 7504 5583
rect 7538 5549 7680 5583
rect 7498 5511 7680 5549
rect 7498 5477 7504 5511
rect 7538 5477 7680 5511
rect 7498 5439 7680 5477
rect 7498 5405 7504 5439
rect 7538 5405 7680 5439
rect 7498 5367 7680 5405
rect 7498 5333 7504 5367
rect 7538 5333 7680 5367
rect 7498 5295 7680 5333
rect 7498 5261 7504 5295
rect 7538 5261 7680 5295
rect 7498 5223 7680 5261
rect 7498 5189 7504 5223
rect 7538 5189 7680 5223
rect 7498 5151 7680 5189
rect 7498 5117 7504 5151
rect 7538 5117 7680 5151
rect 7498 5079 7680 5117
rect 7498 5045 7504 5079
rect 7538 5045 7680 5079
rect 7498 5007 7680 5045
rect 7498 4973 7504 5007
rect 7538 4973 7680 5007
rect 7498 4935 7680 4973
rect 7498 4901 7504 4935
rect 7538 4901 7680 4935
rect 7498 4863 7680 4901
rect 7498 4829 7504 4863
rect 7538 4829 7680 4863
rect 7498 4791 7680 4829
rect 7498 4757 7504 4791
rect 7538 4757 7680 4791
rect 7498 4719 7680 4757
rect 7498 4685 7504 4719
rect 7538 4685 7680 4719
rect 7498 4647 7680 4685
rect 7498 4613 7504 4647
rect 7538 4613 7680 4647
rect 7498 4575 7680 4613
rect 7498 4541 7504 4575
rect 7538 4541 7680 4575
rect 7498 4503 7680 4541
rect 7498 4469 7504 4503
rect 7538 4469 7680 4503
rect 7498 4431 7680 4469
rect 7498 4397 7504 4431
rect 7538 4397 7680 4431
rect 7498 4359 7680 4397
rect 7498 4325 7504 4359
rect 7538 4325 7680 4359
rect 7498 4287 7680 4325
rect 7498 4253 7504 4287
rect 7538 4253 7680 4287
rect 7498 4215 7680 4253
rect 7498 4181 7504 4215
rect 7538 4181 7680 4215
rect 7498 4143 7680 4181
rect 7498 4109 7504 4143
rect 7538 4109 7680 4143
rect 7498 4071 7680 4109
rect 7498 4037 7504 4071
rect 7538 4037 7680 4071
rect 7498 3999 7680 4037
rect 7498 3965 7504 3999
rect 7538 3965 7680 3999
rect 7498 3927 7680 3965
rect 7498 3893 7504 3927
rect 7538 3893 7680 3927
rect 7498 3855 7680 3893
rect 7498 3821 7504 3855
rect 7538 3821 7680 3855
rect 7498 3783 7680 3821
rect 7498 3749 7504 3783
rect 7538 3749 7680 3783
rect 7498 3711 7680 3749
rect 7498 3677 7504 3711
rect 7538 3677 7680 3711
rect 7498 3630 7680 3677
rect 7804 5583 7986 5630
rect 7804 5549 7946 5583
rect 7980 5549 7986 5583
rect 7804 5511 7986 5549
rect 7804 5477 7946 5511
rect 7980 5477 7986 5511
rect 7804 5439 7986 5477
rect 7804 5405 7946 5439
rect 7980 5405 7986 5439
rect 7804 5367 7986 5405
rect 7804 5333 7946 5367
rect 7980 5333 7986 5367
rect 7804 5295 7986 5333
rect 7804 5261 7946 5295
rect 7980 5261 7986 5295
rect 7804 5223 7986 5261
rect 7804 5189 7946 5223
rect 7980 5189 7986 5223
rect 7804 5151 7986 5189
rect 7804 5117 7946 5151
rect 7980 5117 7986 5151
rect 7804 5079 7986 5117
rect 7804 5045 7946 5079
rect 7980 5045 7986 5079
rect 7804 5007 7986 5045
rect 7804 4973 7946 5007
rect 7980 4973 7986 5007
rect 7804 4935 7986 4973
rect 7804 4901 7946 4935
rect 7980 4901 7986 4935
rect 7804 4863 7986 4901
rect 7804 4829 7946 4863
rect 7980 4829 7986 4863
rect 7804 4791 7986 4829
rect 7804 4757 7946 4791
rect 7980 4757 7986 4791
rect 7804 4719 7986 4757
rect 7804 4685 7946 4719
rect 7980 4685 7986 4719
rect 7804 4647 7986 4685
rect 7804 4613 7946 4647
rect 7980 4613 7986 4647
rect 7804 4575 7986 4613
rect 7804 4541 7946 4575
rect 7980 4541 7986 4575
rect 7804 4503 7986 4541
rect 7804 4469 7946 4503
rect 7980 4469 7986 4503
rect 7804 4431 7986 4469
rect 7804 4397 7946 4431
rect 7980 4397 7986 4431
rect 7804 4359 7986 4397
rect 7804 4325 7946 4359
rect 7980 4325 7986 4359
rect 7804 4287 7986 4325
rect 7804 4253 7946 4287
rect 7980 4253 7986 4287
rect 7804 4215 7986 4253
rect 7804 4181 7946 4215
rect 7980 4181 7986 4215
rect 7804 4143 7986 4181
rect 7804 4109 7946 4143
rect 7980 4109 7986 4143
rect 7804 4071 7986 4109
rect 7804 4037 7946 4071
rect 7980 4037 7986 4071
rect 7804 3999 7986 4037
rect 7804 3965 7946 3999
rect 7980 3965 7986 3999
rect 7804 3927 7986 3965
rect 7804 3893 7946 3927
rect 7980 3893 7986 3927
rect 7804 3855 7986 3893
rect 7804 3821 7946 3855
rect 7980 3821 7986 3855
rect 7804 3783 7986 3821
rect 7804 3749 7946 3783
rect 7980 3749 7986 3783
rect 7804 3711 7986 3749
rect 7804 3677 7946 3711
rect 7980 3677 7986 3711
rect 7804 3630 7986 3677
rect 8198 5583 8380 5630
rect 8198 5549 8204 5583
rect 8238 5549 8380 5583
rect 8198 5511 8380 5549
rect 8198 5477 8204 5511
rect 8238 5477 8380 5511
rect 8198 5439 8380 5477
rect 8198 5405 8204 5439
rect 8238 5405 8380 5439
rect 8198 5367 8380 5405
rect 8198 5333 8204 5367
rect 8238 5333 8380 5367
rect 8198 5295 8380 5333
rect 8198 5261 8204 5295
rect 8238 5261 8380 5295
rect 8198 5223 8380 5261
rect 8198 5189 8204 5223
rect 8238 5189 8380 5223
rect 8198 5151 8380 5189
rect 8198 5117 8204 5151
rect 8238 5117 8380 5151
rect 8198 5079 8380 5117
rect 8198 5045 8204 5079
rect 8238 5045 8380 5079
rect 8198 5007 8380 5045
rect 8198 4973 8204 5007
rect 8238 4973 8380 5007
rect 8198 4935 8380 4973
rect 8198 4901 8204 4935
rect 8238 4901 8380 4935
rect 8198 4863 8380 4901
rect 8198 4829 8204 4863
rect 8238 4829 8380 4863
rect 8198 4791 8380 4829
rect 8198 4757 8204 4791
rect 8238 4757 8380 4791
rect 8198 4719 8380 4757
rect 8198 4685 8204 4719
rect 8238 4685 8380 4719
rect 8198 4647 8380 4685
rect 8198 4613 8204 4647
rect 8238 4613 8380 4647
rect 8198 4575 8380 4613
rect 8198 4541 8204 4575
rect 8238 4541 8380 4575
rect 8198 4503 8380 4541
rect 8198 4469 8204 4503
rect 8238 4469 8380 4503
rect 8198 4431 8380 4469
rect 8198 4397 8204 4431
rect 8238 4397 8380 4431
rect 8198 4359 8380 4397
rect 8198 4325 8204 4359
rect 8238 4325 8380 4359
rect 8198 4287 8380 4325
rect 8198 4253 8204 4287
rect 8238 4253 8380 4287
rect 8198 4215 8380 4253
rect 8198 4181 8204 4215
rect 8238 4181 8380 4215
rect 8198 4143 8380 4181
rect 8198 4109 8204 4143
rect 8238 4109 8380 4143
rect 8198 4071 8380 4109
rect 8198 4037 8204 4071
rect 8238 4037 8380 4071
rect 8198 3999 8380 4037
rect 8198 3965 8204 3999
rect 8238 3965 8380 3999
rect 8198 3927 8380 3965
rect 8198 3893 8204 3927
rect 8238 3893 8380 3927
rect 8198 3855 8380 3893
rect 8198 3821 8204 3855
rect 8238 3821 8380 3855
rect 8198 3783 8380 3821
rect 8198 3749 8204 3783
rect 8238 3749 8380 3783
rect 8198 3711 8380 3749
rect 8198 3677 8204 3711
rect 8238 3677 8380 3711
rect 8198 3630 8380 3677
rect 8504 5583 8686 5630
rect 8504 5549 8646 5583
rect 8680 5549 8686 5583
rect 8504 5511 8686 5549
rect 8504 5477 8646 5511
rect 8680 5477 8686 5511
rect 8504 5439 8686 5477
rect 8504 5405 8646 5439
rect 8680 5405 8686 5439
rect 8504 5367 8686 5405
rect 8504 5333 8646 5367
rect 8680 5333 8686 5367
rect 8504 5295 8686 5333
rect 8504 5261 8646 5295
rect 8680 5261 8686 5295
rect 8504 5223 8686 5261
rect 8504 5189 8646 5223
rect 8680 5189 8686 5223
rect 8504 5151 8686 5189
rect 8504 5117 8646 5151
rect 8680 5117 8686 5151
rect 8504 5079 8686 5117
rect 8504 5045 8646 5079
rect 8680 5045 8686 5079
rect 8504 5007 8686 5045
rect 8504 4973 8646 5007
rect 8680 4973 8686 5007
rect 8504 4935 8686 4973
rect 8504 4901 8646 4935
rect 8680 4901 8686 4935
rect 8504 4863 8686 4901
rect 8504 4829 8646 4863
rect 8680 4829 8686 4863
rect 8504 4791 8686 4829
rect 8504 4757 8646 4791
rect 8680 4757 8686 4791
rect 8504 4719 8686 4757
rect 8504 4685 8646 4719
rect 8680 4685 8686 4719
rect 8504 4647 8686 4685
rect 8504 4613 8646 4647
rect 8680 4613 8686 4647
rect 8504 4575 8686 4613
rect 8504 4541 8646 4575
rect 8680 4541 8686 4575
rect 8504 4503 8686 4541
rect 8504 4469 8646 4503
rect 8680 4469 8686 4503
rect 8504 4431 8686 4469
rect 8504 4397 8646 4431
rect 8680 4397 8686 4431
rect 8504 4359 8686 4397
rect 8504 4325 8646 4359
rect 8680 4325 8686 4359
rect 8504 4287 8686 4325
rect 8504 4253 8646 4287
rect 8680 4253 8686 4287
rect 8504 4215 8686 4253
rect 8504 4181 8646 4215
rect 8680 4181 8686 4215
rect 8504 4143 8686 4181
rect 8504 4109 8646 4143
rect 8680 4109 8686 4143
rect 8504 4071 8686 4109
rect 8504 4037 8646 4071
rect 8680 4037 8686 4071
rect 8504 3999 8686 4037
rect 8504 3965 8646 3999
rect 8680 3965 8686 3999
rect 8504 3927 8686 3965
rect 8504 3893 8646 3927
rect 8680 3893 8686 3927
rect 8504 3855 8686 3893
rect 8504 3821 8646 3855
rect 8680 3821 8686 3855
rect 8504 3783 8686 3821
rect 8504 3749 8646 3783
rect 8680 3749 8686 3783
rect 8504 3711 8686 3749
rect 8504 3677 8646 3711
rect 8680 3677 8686 3711
rect 8504 3630 8686 3677
rect 8898 5583 9080 5630
rect 8898 5549 8904 5583
rect 8938 5549 9080 5583
rect 8898 5511 9080 5549
rect 8898 5477 8904 5511
rect 8938 5477 9080 5511
rect 8898 5439 9080 5477
rect 8898 5405 8904 5439
rect 8938 5405 9080 5439
rect 8898 5367 9080 5405
rect 8898 5333 8904 5367
rect 8938 5333 9080 5367
rect 8898 5295 9080 5333
rect 8898 5261 8904 5295
rect 8938 5261 9080 5295
rect 8898 5223 9080 5261
rect 8898 5189 8904 5223
rect 8938 5189 9080 5223
rect 8898 5151 9080 5189
rect 8898 5117 8904 5151
rect 8938 5117 9080 5151
rect 8898 5079 9080 5117
rect 8898 5045 8904 5079
rect 8938 5045 9080 5079
rect 8898 5007 9080 5045
rect 8898 4973 8904 5007
rect 8938 4973 9080 5007
rect 8898 4935 9080 4973
rect 8898 4901 8904 4935
rect 8938 4901 9080 4935
rect 8898 4863 9080 4901
rect 8898 4829 8904 4863
rect 8938 4829 9080 4863
rect 8898 4791 9080 4829
rect 8898 4757 8904 4791
rect 8938 4757 9080 4791
rect 8898 4719 9080 4757
rect 8898 4685 8904 4719
rect 8938 4685 9080 4719
rect 8898 4647 9080 4685
rect 8898 4613 8904 4647
rect 8938 4613 9080 4647
rect 8898 4575 9080 4613
rect 8898 4541 8904 4575
rect 8938 4541 9080 4575
rect 8898 4503 9080 4541
rect 8898 4469 8904 4503
rect 8938 4469 9080 4503
rect 8898 4431 9080 4469
rect 8898 4397 8904 4431
rect 8938 4397 9080 4431
rect 8898 4359 9080 4397
rect 8898 4325 8904 4359
rect 8938 4325 9080 4359
rect 8898 4287 9080 4325
rect 8898 4253 8904 4287
rect 8938 4253 9080 4287
rect 8898 4215 9080 4253
rect 8898 4181 8904 4215
rect 8938 4181 9080 4215
rect 8898 4143 9080 4181
rect 8898 4109 8904 4143
rect 8938 4109 9080 4143
rect 8898 4071 9080 4109
rect 8898 4037 8904 4071
rect 8938 4037 9080 4071
rect 8898 3999 9080 4037
rect 8898 3965 8904 3999
rect 8938 3965 9080 3999
rect 8898 3927 9080 3965
rect 8898 3893 8904 3927
rect 8938 3893 9080 3927
rect 8898 3855 9080 3893
rect 8898 3821 8904 3855
rect 8938 3821 9080 3855
rect 8898 3783 9080 3821
rect 8898 3749 8904 3783
rect 8938 3749 9080 3783
rect 8898 3711 9080 3749
rect 8898 3677 8904 3711
rect 8938 3677 9080 3711
rect 8898 3630 9080 3677
rect 9204 5583 9386 5630
rect 9204 5549 9346 5583
rect 9380 5549 9386 5583
rect 9204 5511 9386 5549
rect 9204 5477 9346 5511
rect 9380 5477 9386 5511
rect 9204 5439 9386 5477
rect 9204 5405 9346 5439
rect 9380 5405 9386 5439
rect 9204 5367 9386 5405
rect 9204 5333 9346 5367
rect 9380 5333 9386 5367
rect 9204 5295 9386 5333
rect 9204 5261 9346 5295
rect 9380 5261 9386 5295
rect 9204 5223 9386 5261
rect 9204 5189 9346 5223
rect 9380 5189 9386 5223
rect 9204 5151 9386 5189
rect 9204 5117 9346 5151
rect 9380 5117 9386 5151
rect 9204 5079 9386 5117
rect 9204 5045 9346 5079
rect 9380 5045 9386 5079
rect 9204 5007 9386 5045
rect 9204 4973 9346 5007
rect 9380 4973 9386 5007
rect 9204 4935 9386 4973
rect 9204 4901 9346 4935
rect 9380 4901 9386 4935
rect 9204 4863 9386 4901
rect 9204 4829 9346 4863
rect 9380 4829 9386 4863
rect 9204 4791 9386 4829
rect 9204 4757 9346 4791
rect 9380 4757 9386 4791
rect 9204 4719 9386 4757
rect 9204 4685 9346 4719
rect 9380 4685 9386 4719
rect 9204 4647 9386 4685
rect 9204 4613 9346 4647
rect 9380 4613 9386 4647
rect 9204 4575 9386 4613
rect 9204 4541 9346 4575
rect 9380 4541 9386 4575
rect 9204 4503 9386 4541
rect 9204 4469 9346 4503
rect 9380 4469 9386 4503
rect 9204 4431 9386 4469
rect 9204 4397 9346 4431
rect 9380 4397 9386 4431
rect 9204 4359 9386 4397
rect 9204 4325 9346 4359
rect 9380 4325 9386 4359
rect 9204 4287 9386 4325
rect 9204 4253 9346 4287
rect 9380 4253 9386 4287
rect 9204 4215 9386 4253
rect 9204 4181 9346 4215
rect 9380 4181 9386 4215
rect 9204 4143 9386 4181
rect 9204 4109 9346 4143
rect 9380 4109 9386 4143
rect 9204 4071 9386 4109
rect 9204 4037 9346 4071
rect 9380 4037 9386 4071
rect 9204 3999 9386 4037
rect 9204 3965 9346 3999
rect 9380 3965 9386 3999
rect 9204 3927 9386 3965
rect 9204 3893 9346 3927
rect 9380 3893 9386 3927
rect 9204 3855 9386 3893
rect 9204 3821 9346 3855
rect 9380 3821 9386 3855
rect 9204 3783 9386 3821
rect 9204 3749 9346 3783
rect 9380 3749 9386 3783
rect 9204 3711 9386 3749
rect 9204 3677 9346 3711
rect 9380 3677 9386 3711
rect 9204 3630 9386 3677
rect 9598 5583 9780 5630
rect 9598 5549 9604 5583
rect 9638 5549 9780 5583
rect 9598 5511 9780 5549
rect 9598 5477 9604 5511
rect 9638 5477 9780 5511
rect 9598 5439 9780 5477
rect 9598 5405 9604 5439
rect 9638 5405 9780 5439
rect 9598 5367 9780 5405
rect 9598 5333 9604 5367
rect 9638 5333 9780 5367
rect 9598 5295 9780 5333
rect 9598 5261 9604 5295
rect 9638 5261 9780 5295
rect 9598 5223 9780 5261
rect 9598 5189 9604 5223
rect 9638 5189 9780 5223
rect 9598 5151 9780 5189
rect 9598 5117 9604 5151
rect 9638 5117 9780 5151
rect 9598 5079 9780 5117
rect 9598 5045 9604 5079
rect 9638 5045 9780 5079
rect 9598 5007 9780 5045
rect 9598 4973 9604 5007
rect 9638 4973 9780 5007
rect 9598 4935 9780 4973
rect 9598 4901 9604 4935
rect 9638 4901 9780 4935
rect 9598 4863 9780 4901
rect 9598 4829 9604 4863
rect 9638 4829 9780 4863
rect 9598 4791 9780 4829
rect 9598 4757 9604 4791
rect 9638 4757 9780 4791
rect 9598 4719 9780 4757
rect 9598 4685 9604 4719
rect 9638 4685 9780 4719
rect 9598 4647 9780 4685
rect 9598 4613 9604 4647
rect 9638 4613 9780 4647
rect 9598 4575 9780 4613
rect 9598 4541 9604 4575
rect 9638 4541 9780 4575
rect 9598 4503 9780 4541
rect 9598 4469 9604 4503
rect 9638 4469 9780 4503
rect 9598 4431 9780 4469
rect 9598 4397 9604 4431
rect 9638 4397 9780 4431
rect 9598 4359 9780 4397
rect 9598 4325 9604 4359
rect 9638 4325 9780 4359
rect 9598 4287 9780 4325
rect 9598 4253 9604 4287
rect 9638 4253 9780 4287
rect 9598 4215 9780 4253
rect 9598 4181 9604 4215
rect 9638 4181 9780 4215
rect 9598 4143 9780 4181
rect 9598 4109 9604 4143
rect 9638 4109 9780 4143
rect 9598 4071 9780 4109
rect 9598 4037 9604 4071
rect 9638 4037 9780 4071
rect 9598 3999 9780 4037
rect 9598 3965 9604 3999
rect 9638 3965 9780 3999
rect 9598 3927 9780 3965
rect 9598 3893 9604 3927
rect 9638 3893 9780 3927
rect 9598 3855 9780 3893
rect 9598 3821 9604 3855
rect 9638 3821 9780 3855
rect 9598 3783 9780 3821
rect 9598 3749 9604 3783
rect 9638 3749 9780 3783
rect 9598 3711 9780 3749
rect 9598 3677 9604 3711
rect 9638 3677 9780 3711
rect 9598 3630 9780 3677
rect 9904 5583 10086 5630
rect 9904 5549 10046 5583
rect 10080 5549 10086 5583
rect 9904 5511 10086 5549
rect 9904 5477 10046 5511
rect 10080 5477 10086 5511
rect 9904 5439 10086 5477
rect 9904 5405 10046 5439
rect 10080 5405 10086 5439
rect 9904 5367 10086 5405
rect 9904 5333 10046 5367
rect 10080 5333 10086 5367
rect 9904 5295 10086 5333
rect 9904 5261 10046 5295
rect 10080 5261 10086 5295
rect 9904 5223 10086 5261
rect 9904 5189 10046 5223
rect 10080 5189 10086 5223
rect 9904 5151 10086 5189
rect 9904 5117 10046 5151
rect 10080 5117 10086 5151
rect 9904 5079 10086 5117
rect 9904 5045 10046 5079
rect 10080 5045 10086 5079
rect 9904 5007 10086 5045
rect 9904 4973 10046 5007
rect 10080 4973 10086 5007
rect 9904 4935 10086 4973
rect 9904 4901 10046 4935
rect 10080 4901 10086 4935
rect 9904 4863 10086 4901
rect 9904 4829 10046 4863
rect 10080 4829 10086 4863
rect 9904 4791 10086 4829
rect 9904 4757 10046 4791
rect 10080 4757 10086 4791
rect 9904 4719 10086 4757
rect 9904 4685 10046 4719
rect 10080 4685 10086 4719
rect 9904 4647 10086 4685
rect 9904 4613 10046 4647
rect 10080 4613 10086 4647
rect 9904 4575 10086 4613
rect 9904 4541 10046 4575
rect 10080 4541 10086 4575
rect 9904 4503 10086 4541
rect 9904 4469 10046 4503
rect 10080 4469 10086 4503
rect 9904 4431 10086 4469
rect 9904 4397 10046 4431
rect 10080 4397 10086 4431
rect 9904 4359 10086 4397
rect 9904 4325 10046 4359
rect 10080 4325 10086 4359
rect 9904 4287 10086 4325
rect 9904 4253 10046 4287
rect 10080 4253 10086 4287
rect 9904 4215 10086 4253
rect 9904 4181 10046 4215
rect 10080 4181 10086 4215
rect 9904 4143 10086 4181
rect 9904 4109 10046 4143
rect 10080 4109 10086 4143
rect 9904 4071 10086 4109
rect 9904 4037 10046 4071
rect 10080 4037 10086 4071
rect 9904 3999 10086 4037
rect 9904 3965 10046 3999
rect 10080 3965 10086 3999
rect 9904 3927 10086 3965
rect 9904 3893 10046 3927
rect 10080 3893 10086 3927
rect 9904 3855 10086 3893
rect 9904 3821 10046 3855
rect 10080 3821 10086 3855
rect 9904 3783 10086 3821
rect 9904 3749 10046 3783
rect 10080 3749 10086 3783
rect 9904 3711 10086 3749
rect 9904 3677 10046 3711
rect 10080 3677 10086 3711
rect 9904 3630 10086 3677
rect 10298 5583 10480 5630
rect 10298 5549 10304 5583
rect 10338 5549 10480 5583
rect 10298 5511 10480 5549
rect 10298 5477 10304 5511
rect 10338 5477 10480 5511
rect 10298 5439 10480 5477
rect 10298 5405 10304 5439
rect 10338 5405 10480 5439
rect 11557 5524 11690 5709
rect 11746 5662 12138 5668
rect 11746 5628 11781 5662
rect 11815 5628 11853 5662
rect 11887 5628 11925 5662
rect 11959 5628 11997 5662
rect 12031 5628 12069 5662
rect 12103 5628 12138 5662
rect 11746 5622 12138 5628
rect 11557 5489 12018 5524
rect 11557 5455 11882 5489
rect 11916 5455 11954 5489
rect 11988 5455 12018 5489
rect 11557 5420 12018 5455
rect 10298 5367 10480 5405
rect 10298 5333 10304 5367
rect 10338 5333 10480 5367
rect 10298 5295 10480 5333
rect 10298 5261 10304 5295
rect 10338 5261 10480 5295
rect 10298 5223 10480 5261
rect 10298 5189 10304 5223
rect 10338 5189 10480 5223
rect 10298 5151 10480 5189
rect 10298 5117 10304 5151
rect 10338 5117 10480 5151
rect 10298 5079 10480 5117
rect 10298 5045 10304 5079
rect 10338 5045 10480 5079
rect 12194 5250 12327 5709
rect 12457 6849 12590 7025
rect 12646 6930 13038 6936
rect 12646 6896 12681 6930
rect 12715 6896 12753 6930
rect 12787 6896 12825 6930
rect 12859 6896 12897 6930
rect 12931 6896 12969 6930
rect 13003 6896 13038 6930
rect 12646 6890 13038 6896
rect 13094 6849 13227 6980
rect 12457 6810 12636 6849
rect 12457 6776 12596 6810
rect 12630 6776 12636 6810
rect 12457 6738 12636 6776
rect 12457 6704 12596 6738
rect 12630 6704 12636 6738
rect 12457 6666 12636 6704
rect 12457 6632 12596 6666
rect 12630 6632 12636 6666
rect 12457 6594 12636 6632
rect 12457 6560 12596 6594
rect 12630 6560 12636 6594
rect 12457 6522 12636 6560
rect 12457 6488 12596 6522
rect 12630 6488 12636 6522
rect 12457 6449 12636 6488
rect 13048 6810 13227 6849
rect 13048 6776 13054 6810
rect 13088 6776 13227 6810
rect 13048 6738 13227 6776
rect 13048 6704 13054 6738
rect 13088 6704 13227 6738
rect 13048 6666 13227 6704
rect 13048 6632 13054 6666
rect 13088 6632 13227 6666
rect 13048 6594 13227 6632
rect 13048 6560 13054 6594
rect 13088 6560 13227 6594
rect 13048 6522 13227 6560
rect 13048 6488 13054 6522
rect 13088 6488 13227 6522
rect 13048 6449 13227 6488
rect 12457 6109 12590 6449
rect 12646 6402 13038 6408
rect 12646 6368 12681 6402
rect 12715 6368 12753 6402
rect 12787 6368 12825 6402
rect 12859 6368 12897 6402
rect 12931 6368 12969 6402
rect 13003 6368 13038 6402
rect 12646 6305 13038 6368
rect 12646 6253 12794 6305
rect 12846 6253 12858 6305
rect 12910 6253 13038 6305
rect 12646 6190 13038 6253
rect 12646 6156 12681 6190
rect 12715 6156 12753 6190
rect 12787 6156 12825 6190
rect 12859 6156 12897 6190
rect 12931 6156 12969 6190
rect 13003 6156 13038 6190
rect 12646 6150 13038 6156
rect 13094 6109 13227 6449
rect 12457 6070 12636 6109
rect 12457 6036 12596 6070
rect 12630 6036 12636 6070
rect 12457 5998 12636 6036
rect 12457 5964 12596 5998
rect 12630 5964 12636 5998
rect 12457 5926 12636 5964
rect 12457 5892 12596 5926
rect 12630 5892 12636 5926
rect 12457 5854 12636 5892
rect 12457 5820 12596 5854
rect 12630 5820 12636 5854
rect 12457 5782 12636 5820
rect 12457 5748 12596 5782
rect 12630 5748 12636 5782
rect 12457 5709 12636 5748
rect 13048 6070 13227 6109
rect 13048 6036 13054 6070
rect 13088 6036 13227 6070
rect 13048 5998 13227 6036
rect 13048 5964 13054 5998
rect 13088 5964 13227 5998
rect 13048 5926 13227 5964
rect 13048 5892 13054 5926
rect 13088 5892 13227 5926
rect 13048 5854 13227 5892
rect 13048 5820 13054 5854
rect 13088 5820 13227 5854
rect 13048 5782 13227 5820
rect 13048 5748 13054 5782
rect 13088 5748 13227 5782
rect 13048 5709 13227 5748
rect 12457 5524 12590 5709
rect 12646 5662 13038 5668
rect 12646 5628 12681 5662
rect 12715 5628 12753 5662
rect 12787 5628 12825 5662
rect 12859 5628 12897 5662
rect 12931 5628 12969 5662
rect 13003 5628 13038 5662
rect 12646 5622 13038 5628
rect 12457 5489 12918 5524
rect 12457 5455 12782 5489
rect 12816 5455 12854 5489
rect 12888 5455 12918 5489
rect 12457 5420 12918 5455
rect 13094 5250 13227 5709
rect 13357 6849 13490 7025
rect 13546 6930 13938 6936
rect 13546 6896 13581 6930
rect 13615 6896 13653 6930
rect 13687 6896 13725 6930
rect 13759 6896 13797 6930
rect 13831 6896 13869 6930
rect 13903 6896 13938 6930
rect 13546 6890 13938 6896
rect 13994 6849 14127 6980
rect 13357 6810 13536 6849
rect 13357 6776 13496 6810
rect 13530 6776 13536 6810
rect 13357 6738 13536 6776
rect 13357 6704 13496 6738
rect 13530 6704 13536 6738
rect 13357 6666 13536 6704
rect 13357 6632 13496 6666
rect 13530 6632 13536 6666
rect 13357 6594 13536 6632
rect 13357 6560 13496 6594
rect 13530 6560 13536 6594
rect 13357 6522 13536 6560
rect 13357 6488 13496 6522
rect 13530 6488 13536 6522
rect 13357 6449 13536 6488
rect 13948 6810 14127 6849
rect 13948 6776 13954 6810
rect 13988 6776 14127 6810
rect 13948 6738 14127 6776
rect 13948 6704 13954 6738
rect 13988 6704 14127 6738
rect 13948 6666 14127 6704
rect 13948 6632 13954 6666
rect 13988 6632 14127 6666
rect 13948 6594 14127 6632
rect 13948 6560 13954 6594
rect 13988 6560 14127 6594
rect 13948 6522 14127 6560
rect 13948 6488 13954 6522
rect 13988 6488 14127 6522
rect 13948 6449 14127 6488
rect 13357 6109 13490 6449
rect 13546 6402 13938 6408
rect 13546 6368 13581 6402
rect 13615 6368 13653 6402
rect 13687 6368 13725 6402
rect 13759 6368 13797 6402
rect 13831 6368 13869 6402
rect 13903 6368 13938 6402
rect 13546 6305 13938 6368
rect 13546 6253 13694 6305
rect 13746 6253 13758 6305
rect 13810 6253 13938 6305
rect 13546 6190 13938 6253
rect 13546 6156 13581 6190
rect 13615 6156 13653 6190
rect 13687 6156 13725 6190
rect 13759 6156 13797 6190
rect 13831 6156 13869 6190
rect 13903 6156 13938 6190
rect 13546 6150 13938 6156
rect 13994 6109 14127 6449
rect 13357 6070 13536 6109
rect 13357 6036 13496 6070
rect 13530 6036 13536 6070
rect 13357 5998 13536 6036
rect 13357 5964 13496 5998
rect 13530 5964 13536 5998
rect 13357 5926 13536 5964
rect 13357 5892 13496 5926
rect 13530 5892 13536 5926
rect 13357 5854 13536 5892
rect 13357 5820 13496 5854
rect 13530 5820 13536 5854
rect 13357 5782 13536 5820
rect 13357 5748 13496 5782
rect 13530 5748 13536 5782
rect 13357 5709 13536 5748
rect 13948 6070 14127 6109
rect 13948 6036 13954 6070
rect 13988 6036 14127 6070
rect 13948 5998 14127 6036
rect 13948 5964 13954 5998
rect 13988 5964 14127 5998
rect 13948 5926 14127 5964
rect 13948 5892 13954 5926
rect 13988 5892 14127 5926
rect 13948 5854 14127 5892
rect 13948 5820 13954 5854
rect 13988 5820 14127 5854
rect 13948 5782 14127 5820
rect 13948 5748 13954 5782
rect 13988 5748 14127 5782
rect 13948 5709 14127 5748
rect 13357 5524 13490 5709
rect 13546 5662 13938 5668
rect 13546 5628 13581 5662
rect 13615 5628 13653 5662
rect 13687 5628 13725 5662
rect 13759 5628 13797 5662
rect 13831 5628 13869 5662
rect 13903 5628 13938 5662
rect 13546 5622 13938 5628
rect 13357 5489 13818 5524
rect 13357 5455 13682 5489
rect 13716 5455 13754 5489
rect 13788 5455 13818 5489
rect 13357 5420 13818 5455
rect 13994 5250 14127 5709
rect 14257 6849 14390 7025
rect 14446 6930 14838 6936
rect 14446 6896 14481 6930
rect 14515 6896 14553 6930
rect 14587 6896 14625 6930
rect 14659 6896 14697 6930
rect 14731 6896 14769 6930
rect 14803 6896 14838 6930
rect 14446 6890 14838 6896
rect 14894 6849 15027 6980
rect 14257 6810 14436 6849
rect 14257 6776 14396 6810
rect 14430 6776 14436 6810
rect 14257 6738 14436 6776
rect 14257 6704 14396 6738
rect 14430 6704 14436 6738
rect 14257 6666 14436 6704
rect 14257 6632 14396 6666
rect 14430 6632 14436 6666
rect 14257 6594 14436 6632
rect 14257 6560 14396 6594
rect 14430 6560 14436 6594
rect 14257 6522 14436 6560
rect 14257 6488 14396 6522
rect 14430 6488 14436 6522
rect 14257 6449 14436 6488
rect 14848 6810 15027 6849
rect 14848 6776 14854 6810
rect 14888 6776 15027 6810
rect 14848 6738 15027 6776
rect 14848 6704 14854 6738
rect 14888 6704 15027 6738
rect 14848 6666 15027 6704
rect 14848 6632 14854 6666
rect 14888 6632 15027 6666
rect 14848 6594 15027 6632
rect 14848 6560 14854 6594
rect 14888 6560 15027 6594
rect 14848 6522 15027 6560
rect 14848 6488 14854 6522
rect 14888 6488 15027 6522
rect 14848 6449 15027 6488
rect 14257 6109 14390 6449
rect 14446 6402 14838 6408
rect 14446 6368 14481 6402
rect 14515 6368 14553 6402
rect 14587 6368 14625 6402
rect 14659 6368 14697 6402
rect 14731 6368 14769 6402
rect 14803 6368 14838 6402
rect 14446 6305 14838 6368
rect 14446 6253 14594 6305
rect 14646 6253 14658 6305
rect 14710 6253 14838 6305
rect 14446 6190 14838 6253
rect 14446 6156 14481 6190
rect 14515 6156 14553 6190
rect 14587 6156 14625 6190
rect 14659 6156 14697 6190
rect 14731 6156 14769 6190
rect 14803 6156 14838 6190
rect 14446 6150 14838 6156
rect 14894 6109 15027 6449
rect 14257 6070 14436 6109
rect 14257 6036 14396 6070
rect 14430 6036 14436 6070
rect 14257 5998 14436 6036
rect 14257 5964 14396 5998
rect 14430 5964 14436 5998
rect 14257 5926 14436 5964
rect 14257 5892 14396 5926
rect 14430 5892 14436 5926
rect 14257 5854 14436 5892
rect 14257 5820 14396 5854
rect 14430 5820 14436 5854
rect 14257 5782 14436 5820
rect 14257 5748 14396 5782
rect 14430 5748 14436 5782
rect 14257 5709 14436 5748
rect 14848 6070 15027 6109
rect 14848 6036 14854 6070
rect 14888 6036 15027 6070
rect 14848 5998 15027 6036
rect 14848 5964 14854 5998
rect 14888 5964 15027 5998
rect 14848 5926 15027 5964
rect 14848 5892 14854 5926
rect 14888 5892 15027 5926
rect 14848 5854 15027 5892
rect 14848 5820 14854 5854
rect 14888 5820 15027 5854
rect 14848 5782 15027 5820
rect 14848 5748 14854 5782
rect 14888 5748 15027 5782
rect 14848 5709 15027 5748
rect 14257 5524 14390 5709
rect 14446 5662 14838 5668
rect 14446 5628 14481 5662
rect 14515 5628 14553 5662
rect 14587 5628 14625 5662
rect 14659 5628 14697 5662
rect 14731 5628 14769 5662
rect 14803 5628 14838 5662
rect 14446 5622 14838 5628
rect 14257 5489 14718 5524
rect 14257 5455 14582 5489
rect 14616 5455 14654 5489
rect 14688 5455 14718 5489
rect 14257 5420 14718 5455
rect 14894 5250 15027 5709
rect 15157 6849 15290 7025
rect 15346 6930 15738 6936
rect 15346 6896 15381 6930
rect 15415 6896 15453 6930
rect 15487 6896 15525 6930
rect 15559 6896 15597 6930
rect 15631 6896 15669 6930
rect 15703 6896 15738 6930
rect 15346 6890 15738 6896
rect 15794 6849 15927 6980
rect 15157 6810 15336 6849
rect 15157 6776 15296 6810
rect 15330 6776 15336 6810
rect 15157 6738 15336 6776
rect 15157 6704 15296 6738
rect 15330 6704 15336 6738
rect 15157 6666 15336 6704
rect 15157 6632 15296 6666
rect 15330 6632 15336 6666
rect 15157 6594 15336 6632
rect 15157 6560 15296 6594
rect 15330 6560 15336 6594
rect 15157 6522 15336 6560
rect 15157 6488 15296 6522
rect 15330 6488 15336 6522
rect 15157 6449 15336 6488
rect 15748 6810 15927 6849
rect 15748 6776 15754 6810
rect 15788 6776 15927 6810
rect 15748 6738 15927 6776
rect 15748 6704 15754 6738
rect 15788 6704 15927 6738
rect 15748 6666 15927 6704
rect 15748 6632 15754 6666
rect 15788 6632 15927 6666
rect 15748 6594 15927 6632
rect 15748 6560 15754 6594
rect 15788 6560 15927 6594
rect 15748 6522 15927 6560
rect 15748 6488 15754 6522
rect 15788 6488 15927 6522
rect 15748 6449 15927 6488
rect 15157 6109 15290 6449
rect 15346 6402 15738 6408
rect 15346 6368 15381 6402
rect 15415 6368 15453 6402
rect 15487 6368 15525 6402
rect 15559 6368 15597 6402
rect 15631 6368 15669 6402
rect 15703 6368 15738 6402
rect 15346 6305 15738 6368
rect 15346 6253 15494 6305
rect 15546 6253 15558 6305
rect 15610 6253 15738 6305
rect 15346 6190 15738 6253
rect 15346 6156 15381 6190
rect 15415 6156 15453 6190
rect 15487 6156 15525 6190
rect 15559 6156 15597 6190
rect 15631 6156 15669 6190
rect 15703 6156 15738 6190
rect 15346 6150 15738 6156
rect 15794 6109 15927 6449
rect 15157 6070 15336 6109
rect 15157 6036 15296 6070
rect 15330 6036 15336 6070
rect 15157 5998 15336 6036
rect 15157 5964 15296 5998
rect 15330 5964 15336 5998
rect 15157 5926 15336 5964
rect 15157 5892 15296 5926
rect 15330 5892 15336 5926
rect 15157 5854 15336 5892
rect 15157 5820 15296 5854
rect 15330 5820 15336 5854
rect 15157 5782 15336 5820
rect 15157 5748 15296 5782
rect 15330 5748 15336 5782
rect 15157 5709 15336 5748
rect 15748 6070 15927 6109
rect 15748 6036 15754 6070
rect 15788 6036 15927 6070
rect 15748 5998 15927 6036
rect 15748 5964 15754 5998
rect 15788 5964 15927 5998
rect 15748 5926 15927 5964
rect 15748 5892 15754 5926
rect 15788 5892 15927 5926
rect 15748 5854 15927 5892
rect 15748 5820 15754 5854
rect 15788 5820 15927 5854
rect 15748 5782 15927 5820
rect 15748 5748 15754 5782
rect 15788 5748 15927 5782
rect 15748 5709 15927 5748
rect 15157 5524 15290 5709
rect 15346 5662 15738 5668
rect 15346 5628 15381 5662
rect 15415 5628 15453 5662
rect 15487 5628 15525 5662
rect 15559 5628 15597 5662
rect 15631 5628 15669 5662
rect 15703 5628 15738 5662
rect 15346 5622 15738 5628
rect 15157 5489 15618 5524
rect 15157 5455 15482 5489
rect 15516 5455 15554 5489
rect 15588 5455 15618 5489
rect 15157 5420 15618 5455
rect 15794 5250 15927 5709
rect 16057 6849 16190 7025
rect 16246 6930 16638 6936
rect 16246 6896 16281 6930
rect 16315 6896 16353 6930
rect 16387 6896 16425 6930
rect 16459 6896 16497 6930
rect 16531 6896 16569 6930
rect 16603 6896 16638 6930
rect 16246 6890 16638 6896
rect 16694 6849 16827 6980
rect 16057 6810 16236 6849
rect 16057 6776 16196 6810
rect 16230 6776 16236 6810
rect 16057 6738 16236 6776
rect 16057 6704 16196 6738
rect 16230 6704 16236 6738
rect 16057 6666 16236 6704
rect 16057 6632 16196 6666
rect 16230 6632 16236 6666
rect 16057 6594 16236 6632
rect 16057 6560 16196 6594
rect 16230 6560 16236 6594
rect 16057 6522 16236 6560
rect 16057 6488 16196 6522
rect 16230 6488 16236 6522
rect 16057 6449 16236 6488
rect 16648 6810 16827 6849
rect 16648 6776 16654 6810
rect 16688 6776 16827 6810
rect 16648 6738 16827 6776
rect 16648 6704 16654 6738
rect 16688 6704 16827 6738
rect 16648 6666 16827 6704
rect 16648 6632 16654 6666
rect 16688 6632 16827 6666
rect 16648 6594 16827 6632
rect 16648 6560 16654 6594
rect 16688 6560 16827 6594
rect 16648 6522 16827 6560
rect 16648 6488 16654 6522
rect 16688 6488 16827 6522
rect 16648 6449 16827 6488
rect 16057 6109 16190 6449
rect 16246 6402 16638 6408
rect 16246 6368 16281 6402
rect 16315 6368 16353 6402
rect 16387 6368 16425 6402
rect 16459 6368 16497 6402
rect 16531 6368 16569 6402
rect 16603 6368 16638 6402
rect 16246 6305 16638 6368
rect 16246 6253 16394 6305
rect 16446 6253 16458 6305
rect 16510 6253 16638 6305
rect 16246 6190 16638 6253
rect 16246 6156 16281 6190
rect 16315 6156 16353 6190
rect 16387 6156 16425 6190
rect 16459 6156 16497 6190
rect 16531 6156 16569 6190
rect 16603 6156 16638 6190
rect 16246 6150 16638 6156
rect 16694 6109 16827 6449
rect 16057 6070 16236 6109
rect 16057 6036 16196 6070
rect 16230 6036 16236 6070
rect 16057 5998 16236 6036
rect 16057 5964 16196 5998
rect 16230 5964 16236 5998
rect 16057 5926 16236 5964
rect 16057 5892 16196 5926
rect 16230 5892 16236 5926
rect 16057 5854 16236 5892
rect 16057 5820 16196 5854
rect 16230 5820 16236 5854
rect 16057 5782 16236 5820
rect 16057 5748 16196 5782
rect 16230 5748 16236 5782
rect 16057 5709 16236 5748
rect 16648 6070 16827 6109
rect 16648 6036 16654 6070
rect 16688 6036 16827 6070
rect 16648 5998 16827 6036
rect 16648 5964 16654 5998
rect 16688 5964 16827 5998
rect 16648 5926 16827 5964
rect 16648 5892 16654 5926
rect 16688 5892 16827 5926
rect 16648 5854 16827 5892
rect 16648 5820 16654 5854
rect 16688 5820 16827 5854
rect 16648 5782 16827 5820
rect 16648 5748 16654 5782
rect 16688 5748 16827 5782
rect 16648 5709 16827 5748
rect 16057 5524 16190 5709
rect 16246 5662 16638 5668
rect 16246 5628 16281 5662
rect 16315 5628 16353 5662
rect 16387 5628 16425 5662
rect 16459 5628 16497 5662
rect 16531 5628 16569 5662
rect 16603 5628 16638 5662
rect 16246 5622 16638 5628
rect 16057 5489 16518 5524
rect 16057 5455 16382 5489
rect 16416 5455 16454 5489
rect 16488 5455 16518 5489
rect 16057 5420 16518 5455
rect 16694 5250 16827 5709
rect 16957 6849 17090 7025
rect 17146 6930 17538 6936
rect 17146 6896 17181 6930
rect 17215 6896 17253 6930
rect 17287 6896 17325 6930
rect 17359 6896 17397 6930
rect 17431 6896 17469 6930
rect 17503 6896 17538 6930
rect 17146 6890 17538 6896
rect 17594 6849 17727 6980
rect 16957 6810 17136 6849
rect 16957 6776 17096 6810
rect 17130 6776 17136 6810
rect 16957 6738 17136 6776
rect 16957 6704 17096 6738
rect 17130 6704 17136 6738
rect 16957 6666 17136 6704
rect 16957 6632 17096 6666
rect 17130 6632 17136 6666
rect 16957 6594 17136 6632
rect 16957 6560 17096 6594
rect 17130 6560 17136 6594
rect 16957 6522 17136 6560
rect 16957 6488 17096 6522
rect 17130 6488 17136 6522
rect 16957 6449 17136 6488
rect 17548 6810 17727 6849
rect 17548 6776 17554 6810
rect 17588 6776 17727 6810
rect 17548 6738 17727 6776
rect 17548 6704 17554 6738
rect 17588 6704 17727 6738
rect 17548 6666 17727 6704
rect 17548 6632 17554 6666
rect 17588 6632 17727 6666
rect 17548 6594 17727 6632
rect 17548 6560 17554 6594
rect 17588 6560 17727 6594
rect 17548 6522 17727 6560
rect 17548 6488 17554 6522
rect 17588 6488 17727 6522
rect 17548 6449 17727 6488
rect 16957 6109 17090 6449
rect 17146 6402 17538 6408
rect 17146 6368 17181 6402
rect 17215 6368 17253 6402
rect 17287 6368 17325 6402
rect 17359 6368 17397 6402
rect 17431 6368 17469 6402
rect 17503 6368 17538 6402
rect 17146 6305 17538 6368
rect 17146 6253 17294 6305
rect 17346 6253 17358 6305
rect 17410 6253 17538 6305
rect 17146 6190 17538 6253
rect 17146 6156 17181 6190
rect 17215 6156 17253 6190
rect 17287 6156 17325 6190
rect 17359 6156 17397 6190
rect 17431 6156 17469 6190
rect 17503 6156 17538 6190
rect 17146 6150 17538 6156
rect 17594 6109 17727 6449
rect 16957 6070 17136 6109
rect 16957 6036 17096 6070
rect 17130 6036 17136 6070
rect 16957 5998 17136 6036
rect 16957 5964 17096 5998
rect 17130 5964 17136 5998
rect 16957 5926 17136 5964
rect 16957 5892 17096 5926
rect 17130 5892 17136 5926
rect 16957 5854 17136 5892
rect 16957 5820 17096 5854
rect 17130 5820 17136 5854
rect 16957 5782 17136 5820
rect 16957 5748 17096 5782
rect 17130 5748 17136 5782
rect 16957 5709 17136 5748
rect 17548 6070 17727 6109
rect 17548 6036 17554 6070
rect 17588 6036 17727 6070
rect 17548 5998 17727 6036
rect 17548 5964 17554 5998
rect 17588 5964 17727 5998
rect 17548 5926 17727 5964
rect 17548 5892 17554 5926
rect 17588 5892 17727 5926
rect 17548 5854 17727 5892
rect 17548 5820 17554 5854
rect 17588 5820 17727 5854
rect 17548 5782 17727 5820
rect 17548 5748 17554 5782
rect 17588 5748 17727 5782
rect 17548 5709 17727 5748
rect 16957 5524 17090 5709
rect 17146 5662 17538 5668
rect 17146 5628 17181 5662
rect 17215 5628 17253 5662
rect 17287 5628 17325 5662
rect 17359 5628 17397 5662
rect 17431 5628 17469 5662
rect 17503 5628 17538 5662
rect 17146 5622 17538 5628
rect 16957 5489 17418 5524
rect 16957 5455 17282 5489
rect 17316 5455 17354 5489
rect 17388 5455 17418 5489
rect 16957 5420 17418 5455
rect 17594 5250 17727 5709
rect 17857 6849 17990 7025
rect 18046 6930 18438 6936
rect 18046 6896 18081 6930
rect 18115 6896 18153 6930
rect 18187 6896 18225 6930
rect 18259 6896 18297 6930
rect 18331 6896 18369 6930
rect 18403 6896 18438 6930
rect 18046 6890 18438 6896
rect 18494 6849 18627 6980
rect 17857 6810 18036 6849
rect 17857 6776 17996 6810
rect 18030 6776 18036 6810
rect 17857 6738 18036 6776
rect 17857 6704 17996 6738
rect 18030 6704 18036 6738
rect 17857 6666 18036 6704
rect 17857 6632 17996 6666
rect 18030 6632 18036 6666
rect 17857 6594 18036 6632
rect 17857 6560 17996 6594
rect 18030 6560 18036 6594
rect 17857 6522 18036 6560
rect 17857 6488 17996 6522
rect 18030 6488 18036 6522
rect 17857 6449 18036 6488
rect 18448 6810 18627 6849
rect 18448 6776 18454 6810
rect 18488 6776 18627 6810
rect 18448 6738 18627 6776
rect 18448 6704 18454 6738
rect 18488 6704 18627 6738
rect 18448 6666 18627 6704
rect 18448 6632 18454 6666
rect 18488 6632 18627 6666
rect 18448 6594 18627 6632
rect 18448 6560 18454 6594
rect 18488 6560 18627 6594
rect 18448 6522 18627 6560
rect 18448 6488 18454 6522
rect 18488 6488 18627 6522
rect 18448 6449 18627 6488
rect 17857 6109 17990 6449
rect 18046 6402 18438 6408
rect 18046 6368 18081 6402
rect 18115 6368 18153 6402
rect 18187 6368 18225 6402
rect 18259 6368 18297 6402
rect 18331 6368 18369 6402
rect 18403 6368 18438 6402
rect 18046 6305 18438 6368
rect 18046 6253 18194 6305
rect 18246 6253 18258 6305
rect 18310 6253 18438 6305
rect 18046 6190 18438 6253
rect 18046 6156 18081 6190
rect 18115 6156 18153 6190
rect 18187 6156 18225 6190
rect 18259 6156 18297 6190
rect 18331 6156 18369 6190
rect 18403 6156 18438 6190
rect 18046 6150 18438 6156
rect 18494 6109 18627 6449
rect 17857 6070 18036 6109
rect 17857 6036 17996 6070
rect 18030 6036 18036 6070
rect 17857 5998 18036 6036
rect 17857 5964 17996 5998
rect 18030 5964 18036 5998
rect 17857 5926 18036 5964
rect 17857 5892 17996 5926
rect 18030 5892 18036 5926
rect 17857 5854 18036 5892
rect 17857 5820 17996 5854
rect 18030 5820 18036 5854
rect 17857 5782 18036 5820
rect 17857 5748 17996 5782
rect 18030 5748 18036 5782
rect 17857 5709 18036 5748
rect 18448 6070 18627 6109
rect 18448 6036 18454 6070
rect 18488 6036 18627 6070
rect 18448 5998 18627 6036
rect 18448 5964 18454 5998
rect 18488 5964 18627 5998
rect 18448 5926 18627 5964
rect 18448 5892 18454 5926
rect 18488 5892 18627 5926
rect 18448 5854 18627 5892
rect 18448 5820 18454 5854
rect 18488 5820 18627 5854
rect 21073 5982 21155 7496
rect 21073 5930 21089 5982
rect 21141 5930 21155 5982
rect 21073 5918 21155 5930
rect 21073 5866 21089 5918
rect 21141 5866 21155 5918
rect 21073 5853 21155 5866
rect 21449 6469 21567 6483
rect 21449 6075 21455 6469
rect 21561 6075 21567 6469
rect 18448 5782 18627 5820
rect 18448 5748 18454 5782
rect 18488 5748 18627 5782
rect 18448 5709 18627 5748
rect 17857 5524 17990 5709
rect 18046 5662 18438 5668
rect 18046 5628 18081 5662
rect 18115 5628 18153 5662
rect 18187 5628 18225 5662
rect 18259 5628 18297 5662
rect 18331 5628 18369 5662
rect 18403 5628 18438 5662
rect 18046 5622 18438 5628
rect 17857 5489 18318 5524
rect 17857 5455 18182 5489
rect 18216 5455 18254 5489
rect 18288 5455 18318 5489
rect 17857 5420 18318 5455
rect 18494 5250 18627 5709
rect 12194 5064 18627 5250
rect 10298 5007 10480 5045
rect 10298 4973 10304 5007
rect 10338 4973 10480 5007
rect 10298 4935 10480 4973
rect 10298 4901 10304 4935
rect 10338 4901 10480 4935
rect 10298 4863 10480 4901
rect 10298 4829 10304 4863
rect 10338 4829 10480 4863
rect 10298 4791 10480 4829
rect 10298 4757 10304 4791
rect 10338 4757 10480 4791
rect 10298 4719 10480 4757
rect 10298 4685 10304 4719
rect 10338 4685 10480 4719
rect 10298 4647 10480 4685
rect 10298 4613 10304 4647
rect 10338 4613 10480 4647
rect 10298 4575 10480 4613
rect 10298 4541 10304 4575
rect 10338 4541 10480 4575
rect 10298 4503 10480 4541
rect 10298 4469 10304 4503
rect 10338 4469 10480 4503
rect 10298 4431 10480 4469
rect 10298 4397 10304 4431
rect 10338 4397 10480 4431
rect 10298 4359 10480 4397
rect 10298 4325 10304 4359
rect 10338 4325 10480 4359
rect 10298 4287 10480 4325
rect 10298 4253 10304 4287
rect 10338 4253 10480 4287
rect 10298 4215 10480 4253
rect 10298 4181 10304 4215
rect 10338 4181 10480 4215
rect 10298 4143 10480 4181
rect 10298 4109 10304 4143
rect 10338 4109 10480 4143
rect 10298 4071 10480 4109
rect 10298 4037 10304 4071
rect 10338 4037 10480 4071
rect 10298 3999 10480 4037
rect 10298 3965 10304 3999
rect 10338 3965 10480 3999
rect 10298 3927 10480 3965
rect 10298 3893 10304 3927
rect 10338 3893 10480 3927
rect 10298 3855 10480 3893
rect 10298 3821 10304 3855
rect 10338 3821 10480 3855
rect 10298 3783 10480 3821
rect 10298 3749 10304 3783
rect 10338 3749 10480 3783
rect 10298 3711 10480 3749
rect 10298 3677 10304 3711
rect 10338 3677 10480 3711
rect 10298 3630 10480 3677
rect -4204 3592 -4012 3598
rect -4204 3558 -4161 3592
rect -4127 3558 -4089 3592
rect -4055 3558 -4012 3592
rect -4204 3483 -4012 3558
rect -4204 3431 -4165 3483
rect -4113 3431 -4101 3483
rect -4049 3431 -4012 3483
rect -4204 3357 -4012 3431
rect -3956 3080 -3820 3630
rect -3504 3592 -3312 3598
rect -3504 3558 -3461 3592
rect -3427 3558 -3389 3592
rect -3355 3558 -3312 3592
rect -3504 3483 -3312 3558
rect -3504 3431 -3465 3483
rect -3413 3431 -3401 3483
rect -3349 3431 -3312 3483
rect -3504 3357 -3312 3431
rect -3256 3080 -3120 3630
rect -2804 3592 -2612 3598
rect -2804 3558 -2761 3592
rect -2727 3558 -2689 3592
rect -2655 3558 -2612 3592
rect -2804 3483 -2612 3558
rect -2804 3431 -2765 3483
rect -2713 3431 -2701 3483
rect -2649 3431 -2612 3483
rect -2804 3357 -2612 3431
rect -2556 3080 -2420 3630
rect -2104 3592 -1912 3598
rect -2104 3558 -2061 3592
rect -2027 3558 -1989 3592
rect -1955 3558 -1912 3592
rect -2104 3483 -1912 3558
rect -2104 3431 -2065 3483
rect -2013 3431 -2001 3483
rect -1949 3431 -1912 3483
rect -2104 3357 -1912 3431
rect -1856 3080 -1720 3630
rect -1404 3592 -1212 3598
rect -1404 3558 -1361 3592
rect -1327 3558 -1289 3592
rect -1255 3558 -1212 3592
rect -1404 3483 -1212 3558
rect -1404 3431 -1365 3483
rect -1313 3431 -1301 3483
rect -1249 3431 -1212 3483
rect -1404 3357 -1212 3431
rect -1156 3080 -1020 3630
rect -704 3592 -512 3598
rect -704 3558 -661 3592
rect -627 3558 -589 3592
rect -555 3558 -512 3592
rect -704 3483 -512 3558
rect -704 3431 -665 3483
rect -613 3431 -601 3483
rect -549 3431 -512 3483
rect -704 3357 -512 3431
rect -456 3080 -320 3630
rect -4 3592 188 3598
rect -4 3558 39 3592
rect 73 3558 111 3592
rect 145 3558 188 3592
rect -4 3483 188 3558
rect -4 3431 35 3483
rect 87 3431 99 3483
rect 151 3431 188 3483
rect -4 3357 188 3431
rect 244 3080 380 3630
rect 696 3592 888 3598
rect 696 3558 739 3592
rect 773 3558 811 3592
rect 845 3558 888 3592
rect 696 3483 888 3558
rect 696 3431 735 3483
rect 787 3431 799 3483
rect 851 3431 888 3483
rect 696 3357 888 3431
rect 944 3080 1080 3630
rect 1396 3592 1588 3598
rect 1396 3558 1439 3592
rect 1473 3558 1511 3592
rect 1545 3558 1588 3592
rect 1396 3483 1588 3558
rect 1396 3431 1435 3483
rect 1487 3431 1499 3483
rect 1551 3431 1588 3483
rect 1396 3357 1588 3431
rect 1644 3080 1780 3630
rect 2096 3592 2288 3598
rect 2096 3558 2139 3592
rect 2173 3558 2211 3592
rect 2245 3558 2288 3592
rect 2096 3483 2288 3558
rect 2096 3431 2135 3483
rect 2187 3431 2199 3483
rect 2251 3431 2288 3483
rect 2096 3357 2288 3431
rect 2344 3080 2480 3630
rect 3796 3592 3988 3598
rect 3796 3558 3839 3592
rect 3873 3558 3911 3592
rect 3945 3558 3988 3592
rect 3796 3483 3988 3558
rect 3796 3431 3835 3483
rect 3887 3431 3899 3483
rect 3951 3431 3988 3483
rect 3796 3357 3988 3431
rect 4044 3080 4180 3630
rect 4496 3592 4688 3598
rect 4496 3558 4539 3592
rect 4573 3558 4611 3592
rect 4645 3558 4688 3592
rect 4496 3483 4688 3558
rect 4496 3431 4535 3483
rect 4587 3431 4599 3483
rect 4651 3431 4688 3483
rect 4496 3357 4688 3431
rect 4744 3080 4880 3630
rect 5196 3592 5388 3598
rect 5196 3558 5239 3592
rect 5273 3558 5311 3592
rect 5345 3558 5388 3592
rect 5196 3483 5388 3558
rect 5196 3431 5235 3483
rect 5287 3431 5299 3483
rect 5351 3431 5388 3483
rect 5196 3357 5388 3431
rect 5444 3080 5580 3630
rect 5896 3592 6088 3598
rect 5896 3558 5939 3592
rect 5973 3558 6011 3592
rect 6045 3558 6088 3592
rect 5896 3483 6088 3558
rect 5896 3431 5935 3483
rect 5987 3431 5999 3483
rect 6051 3431 6088 3483
rect 5896 3357 6088 3431
rect 6144 3080 6280 3630
rect 6596 3592 6788 3598
rect 6596 3558 6639 3592
rect 6673 3558 6711 3592
rect 6745 3558 6788 3592
rect 6596 3483 6788 3558
rect 6596 3431 6635 3483
rect 6687 3431 6699 3483
rect 6751 3431 6788 3483
rect 6596 3357 6788 3431
rect 6844 3080 6980 3630
rect 7296 3592 7488 3598
rect 7296 3558 7339 3592
rect 7373 3558 7411 3592
rect 7445 3558 7488 3592
rect 7296 3483 7488 3558
rect 7296 3431 7335 3483
rect 7387 3431 7399 3483
rect 7451 3431 7488 3483
rect 7296 3357 7488 3431
rect 7544 3080 7680 3630
rect 7996 3592 8188 3598
rect 7996 3558 8039 3592
rect 8073 3558 8111 3592
rect 8145 3558 8188 3592
rect 7996 3483 8188 3558
rect 7996 3431 8035 3483
rect 8087 3431 8099 3483
rect 8151 3431 8188 3483
rect 7996 3357 8188 3431
rect 8244 3080 8380 3630
rect 8696 3592 8888 3598
rect 8696 3558 8739 3592
rect 8773 3558 8811 3592
rect 8845 3558 8888 3592
rect 8696 3483 8888 3558
rect 8696 3431 8735 3483
rect 8787 3431 8799 3483
rect 8851 3431 8888 3483
rect 8696 3357 8888 3431
rect 8944 3080 9080 3630
rect 9396 3592 9588 3598
rect 9396 3558 9439 3592
rect 9473 3558 9511 3592
rect 9545 3558 9588 3592
rect 9396 3483 9588 3558
rect 9396 3431 9435 3483
rect 9487 3431 9499 3483
rect 9551 3431 9588 3483
rect 9396 3357 9588 3431
rect 9644 3080 9780 3630
rect 10096 3592 10288 3598
rect 10096 3558 10139 3592
rect 10173 3558 10211 3592
rect 10245 3558 10288 3592
rect 10096 3483 10288 3558
rect 10096 3431 10135 3483
rect 10187 3431 10199 3483
rect 10251 3431 10288 3483
rect 10096 3357 10288 3431
rect 10344 3080 10480 3630
rect -3956 2920 10480 3080
rect 12291 3975 12461 5064
rect 21449 3975 21567 6075
rect 33530 3975 33850 3980
rect 12291 3739 33850 3975
rect -4794 2699 -4767 2751
rect -4715 2699 -4689 2751
rect -4794 2687 -4689 2699
rect -4794 2635 -4767 2687
rect -4715 2635 -4689 2687
rect -4794 2613 -4689 2635
rect -9200 2411 -9070 2420
rect -9200 2287 1711 2411
rect -9200 2280 -9070 2287
rect 1273 2142 1403 2146
rect 957 2134 1403 2142
rect 957 2100 1285 2134
rect 1319 2100 1357 2134
rect 1391 2100 1403 2134
rect 957 2088 1403 2100
rect 957 2075 1401 2088
rect 957 1916 1082 2075
rect 1138 1988 1530 1994
rect 1138 1954 1173 1988
rect 1207 1954 1245 1988
rect 1279 1954 1317 1988
rect 1351 1954 1389 1988
rect 1423 1954 1461 1988
rect 1495 1954 1530 1988
rect 1138 1948 1530 1954
rect 1586 1916 1711 2287
rect 2273 2142 2403 2146
rect 957 1869 1128 1916
rect 957 1835 1088 1869
rect 1122 1835 1128 1869
rect 957 1797 1128 1835
rect 957 1763 1088 1797
rect 1122 1763 1128 1797
rect 957 1716 1128 1763
rect 1540 1869 1711 1916
rect 1540 1835 1546 1869
rect 1580 1835 1711 1869
rect 1540 1797 1711 1835
rect 1540 1763 1546 1797
rect 1580 1763 1711 1797
rect 1540 1716 1711 1763
rect 957 1416 1082 1716
rect 1138 1678 1530 1684
rect 1138 1644 1173 1678
rect 1207 1644 1245 1678
rect 1279 1644 1317 1678
rect 1351 1644 1389 1678
rect 1423 1644 1461 1678
rect 1495 1644 1530 1678
rect 1138 1637 1530 1644
rect 1586 1637 1711 1716
rect 1138 1593 1711 1637
rect 1138 1541 1283 1593
rect 1335 1541 1347 1593
rect 1399 1541 1711 1593
rect 1138 1493 1711 1541
rect 1138 1488 1530 1493
rect 1138 1454 1173 1488
rect 1207 1454 1245 1488
rect 1279 1454 1317 1488
rect 1351 1454 1389 1488
rect 1423 1454 1461 1488
rect 1495 1454 1530 1488
rect 1138 1448 1530 1454
rect 1586 1416 1711 1493
rect 957 1369 1128 1416
rect 957 1335 1088 1369
rect 1122 1335 1128 1369
rect 957 1297 1128 1335
rect 957 1263 1088 1297
rect 1122 1263 1128 1297
rect 957 1216 1128 1263
rect 1540 1369 1711 1416
rect 1540 1335 1546 1369
rect 1580 1335 1711 1369
rect 1540 1297 1711 1335
rect 1540 1263 1546 1297
rect 1580 1263 1711 1297
rect 1540 1216 1711 1263
rect 957 1010 1082 1216
rect 1138 1178 1530 1184
rect 1138 1144 1173 1178
rect 1207 1144 1245 1178
rect 1279 1144 1317 1178
rect 1351 1144 1389 1178
rect 1423 1144 1461 1178
rect 1495 1144 1530 1178
rect 1138 1138 1530 1144
rect 957 1009 1401 1010
rect 957 997 1402 1009
rect 957 963 1284 997
rect 1318 963 1356 997
rect 1390 963 1402 997
rect 957 951 1402 963
rect 957 943 1401 951
rect -9200 713 -8990 720
rect 957 713 1082 943
rect 1586 860 1711 1216
rect 1957 2134 2403 2142
rect 1957 2100 2285 2134
rect 2319 2100 2357 2134
rect 2391 2100 2403 2134
rect 1957 2088 2403 2100
rect 1957 2075 2401 2088
rect 1957 1916 2082 2075
rect 2138 1988 2530 1994
rect 2138 1954 2173 1988
rect 2207 1954 2245 1988
rect 2279 1954 2317 1988
rect 2351 1954 2389 1988
rect 2423 1954 2461 1988
rect 2495 1954 2530 1988
rect 2138 1948 2530 1954
rect 2586 1916 2711 2920
rect 12291 2520 12461 3739
rect 33530 3730 33850 3739
rect 3586 2397 12461 2520
rect 3273 2142 3403 2146
rect 1957 1869 2128 1916
rect 1957 1835 2088 1869
rect 2122 1835 2128 1869
rect 1957 1797 2128 1835
rect 1957 1763 2088 1797
rect 2122 1763 2128 1797
rect 1957 1716 2128 1763
rect 2540 1869 2711 1916
rect 2540 1835 2546 1869
rect 2580 1835 2711 1869
rect 2540 1797 2711 1835
rect 2540 1763 2546 1797
rect 2580 1763 2711 1797
rect 2540 1716 2711 1763
rect 1957 1416 2082 1716
rect 2138 1678 2530 1684
rect 2138 1644 2173 1678
rect 2207 1644 2245 1678
rect 2279 1644 2317 1678
rect 2351 1644 2389 1678
rect 2423 1644 2461 1678
rect 2495 1644 2530 1678
rect 2138 1593 2530 1644
rect 2138 1541 2283 1593
rect 2335 1541 2347 1593
rect 2399 1541 2530 1593
rect 2138 1488 2530 1541
rect 2138 1454 2173 1488
rect 2207 1454 2245 1488
rect 2279 1454 2317 1488
rect 2351 1454 2389 1488
rect 2423 1454 2461 1488
rect 2495 1454 2530 1488
rect 2138 1448 2530 1454
rect 2586 1416 2711 1716
rect 1957 1369 2128 1416
rect 1957 1335 2088 1369
rect 2122 1335 2128 1369
rect 1957 1297 2128 1335
rect 1957 1263 2088 1297
rect 2122 1263 2128 1297
rect 1957 1216 2128 1263
rect 2540 1369 2711 1416
rect 2540 1335 2546 1369
rect 2580 1335 2711 1369
rect 2540 1297 2711 1335
rect 2540 1263 2546 1297
rect 2580 1263 2711 1297
rect 2540 1216 2711 1263
rect 1957 1010 2082 1216
rect 2138 1178 2530 1184
rect 2138 1144 2173 1178
rect 2207 1144 2245 1178
rect 2279 1144 2317 1178
rect 2351 1144 2389 1178
rect 2423 1144 2461 1178
rect 2495 1144 2530 1178
rect 2138 1138 2530 1144
rect 1957 1009 2401 1010
rect 1957 997 2402 1009
rect 1957 963 2284 997
rect 2318 963 2356 997
rect 2390 963 2402 997
rect 1957 951 2402 963
rect 1957 943 2401 951
rect 1957 713 2082 943
rect 2586 860 2711 1216
rect 2957 2134 3403 2142
rect 2957 2100 3285 2134
rect 3319 2100 3357 2134
rect 3391 2100 3403 2134
rect 2957 2088 3403 2100
rect 2957 2075 3401 2088
rect 2957 1916 3082 2075
rect 3138 1988 3530 1994
rect 3138 1954 3173 1988
rect 3207 1954 3245 1988
rect 3279 1954 3317 1988
rect 3351 1954 3389 1988
rect 3423 1954 3461 1988
rect 3495 1954 3530 1988
rect 3138 1948 3530 1954
rect 3586 1916 3711 2397
rect 4273 2142 4403 2146
rect 2957 1869 3128 1916
rect 2957 1835 3088 1869
rect 3122 1835 3128 1869
rect 2957 1797 3128 1835
rect 2957 1763 3088 1797
rect 3122 1763 3128 1797
rect 2957 1716 3128 1763
rect 3540 1869 3711 1916
rect 3540 1835 3546 1869
rect 3580 1835 3711 1869
rect 3540 1797 3711 1835
rect 3540 1763 3546 1797
rect 3580 1763 3711 1797
rect 3540 1716 3711 1763
rect 2957 1416 3082 1716
rect 3138 1678 3530 1684
rect 3138 1644 3173 1678
rect 3207 1644 3245 1678
rect 3279 1644 3317 1678
rect 3351 1644 3389 1678
rect 3423 1644 3461 1678
rect 3495 1644 3530 1678
rect 3138 1593 3530 1644
rect 3138 1541 3283 1593
rect 3335 1541 3347 1593
rect 3399 1541 3530 1593
rect 3138 1488 3530 1541
rect 3138 1454 3173 1488
rect 3207 1454 3245 1488
rect 3279 1454 3317 1488
rect 3351 1454 3389 1488
rect 3423 1454 3461 1488
rect 3495 1454 3530 1488
rect 3138 1448 3530 1454
rect 3586 1416 3711 1716
rect 2957 1369 3128 1416
rect 2957 1335 3088 1369
rect 3122 1335 3128 1369
rect 2957 1297 3128 1335
rect 2957 1263 3088 1297
rect 3122 1263 3128 1297
rect 2957 1216 3128 1263
rect 3540 1369 3711 1416
rect 3540 1335 3546 1369
rect 3580 1335 3711 1369
rect 3540 1297 3711 1335
rect 3540 1263 3546 1297
rect 3580 1263 3711 1297
rect 3540 1216 3711 1263
rect 2957 1010 3082 1216
rect 3138 1178 3530 1184
rect 3138 1144 3173 1178
rect 3207 1144 3245 1178
rect 3279 1144 3317 1178
rect 3351 1144 3389 1178
rect 3423 1144 3461 1178
rect 3495 1144 3530 1178
rect 3138 1138 3530 1144
rect 2957 1009 3401 1010
rect 2957 997 3402 1009
rect 2957 963 3284 997
rect 3318 963 3356 997
rect 3390 963 3402 997
rect 2957 951 3402 963
rect 2957 943 3401 951
rect 2957 713 3082 943
rect 3586 860 3711 1216
rect 3957 2134 4403 2142
rect 3957 2100 4285 2134
rect 4319 2100 4357 2134
rect 4391 2100 4403 2134
rect 3957 2088 4403 2100
rect 3957 2075 4401 2088
rect 3957 1916 4082 2075
rect 4138 1988 4530 1994
rect 4138 1954 4173 1988
rect 4207 1954 4245 1988
rect 4279 1954 4317 1988
rect 4351 1954 4389 1988
rect 4423 1954 4461 1988
rect 4495 1954 4530 1988
rect 4138 1948 4530 1954
rect 4586 1916 4711 2397
rect 5273 2142 5403 2146
rect 3957 1869 4128 1916
rect 3957 1835 4088 1869
rect 4122 1835 4128 1869
rect 3957 1797 4128 1835
rect 3957 1763 4088 1797
rect 4122 1763 4128 1797
rect 3957 1716 4128 1763
rect 4540 1869 4711 1916
rect 4540 1835 4546 1869
rect 4580 1835 4711 1869
rect 4540 1797 4711 1835
rect 4540 1763 4546 1797
rect 4580 1763 4711 1797
rect 4540 1716 4711 1763
rect 3957 1416 4082 1716
rect 4138 1678 4530 1684
rect 4138 1644 4173 1678
rect 4207 1644 4245 1678
rect 4279 1644 4317 1678
rect 4351 1644 4389 1678
rect 4423 1644 4461 1678
rect 4495 1644 4530 1678
rect 4138 1593 4530 1644
rect 4138 1541 4283 1593
rect 4335 1541 4347 1593
rect 4399 1541 4530 1593
rect 4138 1488 4530 1541
rect 4138 1454 4173 1488
rect 4207 1454 4245 1488
rect 4279 1454 4317 1488
rect 4351 1454 4389 1488
rect 4423 1454 4461 1488
rect 4495 1454 4530 1488
rect 4138 1448 4530 1454
rect 4586 1416 4711 1716
rect 3957 1369 4128 1416
rect 3957 1335 4088 1369
rect 4122 1335 4128 1369
rect 3957 1297 4128 1335
rect 3957 1263 4088 1297
rect 4122 1263 4128 1297
rect 3957 1216 4128 1263
rect 4540 1369 4711 1416
rect 4540 1335 4546 1369
rect 4580 1335 4711 1369
rect 4540 1297 4711 1335
rect 4540 1263 4546 1297
rect 4580 1263 4711 1297
rect 4540 1216 4711 1263
rect 3957 1010 4082 1216
rect 4138 1178 4530 1184
rect 4138 1144 4173 1178
rect 4207 1144 4245 1178
rect 4279 1144 4317 1178
rect 4351 1144 4389 1178
rect 4423 1144 4461 1178
rect 4495 1144 4530 1178
rect 4138 1138 4530 1144
rect 3957 1009 4401 1010
rect 3957 997 4402 1009
rect 3957 963 4284 997
rect 4318 963 4356 997
rect 4390 963 4402 997
rect 3957 951 4402 963
rect 3957 943 4401 951
rect 3957 713 4082 943
rect 4586 860 4711 1216
rect 4957 2134 5403 2142
rect 4957 2100 5285 2134
rect 5319 2100 5357 2134
rect 5391 2100 5403 2134
rect 4957 2088 5403 2100
rect 4957 2075 5401 2088
rect 4957 1916 5082 2075
rect 5138 1988 5530 1994
rect 5138 1954 5173 1988
rect 5207 1954 5245 1988
rect 5279 1954 5317 1988
rect 5351 1954 5389 1988
rect 5423 1954 5461 1988
rect 5495 1954 5530 1988
rect 5138 1948 5530 1954
rect 5586 1916 5711 2397
rect 6273 2142 6403 2146
rect 4957 1869 5128 1916
rect 4957 1835 5088 1869
rect 5122 1835 5128 1869
rect 4957 1797 5128 1835
rect 4957 1763 5088 1797
rect 5122 1763 5128 1797
rect 4957 1716 5128 1763
rect 5540 1869 5711 1916
rect 5540 1835 5546 1869
rect 5580 1835 5711 1869
rect 5540 1797 5711 1835
rect 5540 1763 5546 1797
rect 5580 1763 5711 1797
rect 5540 1716 5711 1763
rect 4957 1416 5082 1716
rect 5138 1678 5530 1684
rect 5138 1644 5173 1678
rect 5207 1644 5245 1678
rect 5279 1644 5317 1678
rect 5351 1644 5389 1678
rect 5423 1644 5461 1678
rect 5495 1644 5530 1678
rect 5138 1593 5530 1644
rect 5138 1541 5283 1593
rect 5335 1541 5347 1593
rect 5399 1541 5530 1593
rect 5138 1488 5530 1541
rect 5138 1454 5173 1488
rect 5207 1454 5245 1488
rect 5279 1454 5317 1488
rect 5351 1454 5389 1488
rect 5423 1454 5461 1488
rect 5495 1454 5530 1488
rect 5138 1448 5530 1454
rect 5586 1416 5711 1716
rect 4957 1369 5128 1416
rect 4957 1335 5088 1369
rect 5122 1335 5128 1369
rect 4957 1297 5128 1335
rect 4957 1263 5088 1297
rect 5122 1263 5128 1297
rect 4957 1216 5128 1263
rect 5540 1369 5711 1416
rect 5540 1335 5546 1369
rect 5580 1335 5711 1369
rect 5540 1297 5711 1335
rect 5540 1263 5546 1297
rect 5580 1263 5711 1297
rect 5540 1216 5711 1263
rect 4957 1010 5082 1216
rect 5138 1178 5530 1184
rect 5138 1144 5173 1178
rect 5207 1144 5245 1178
rect 5279 1144 5317 1178
rect 5351 1144 5389 1178
rect 5423 1144 5461 1178
rect 5495 1144 5530 1178
rect 5138 1138 5530 1144
rect 4957 1009 5401 1010
rect 4957 997 5402 1009
rect 4957 963 5284 997
rect 5318 963 5356 997
rect 5390 963 5402 997
rect 4957 951 5402 963
rect 4957 943 5401 951
rect 4957 713 5082 943
rect 5586 860 5711 1216
rect 5957 2134 6403 2142
rect 5957 2100 6285 2134
rect 6319 2100 6357 2134
rect 6391 2100 6403 2134
rect 5957 2088 6403 2100
rect 5957 2075 6401 2088
rect 5957 1916 6082 2075
rect 6138 1988 6530 1994
rect 6138 1954 6173 1988
rect 6207 1954 6245 1988
rect 6279 1954 6317 1988
rect 6351 1954 6389 1988
rect 6423 1954 6461 1988
rect 6495 1954 6530 1988
rect 6138 1948 6530 1954
rect 6586 1916 6711 2397
rect 7273 2142 7403 2146
rect 5957 1869 6128 1916
rect 5957 1835 6088 1869
rect 6122 1835 6128 1869
rect 5957 1797 6128 1835
rect 5957 1763 6088 1797
rect 6122 1763 6128 1797
rect 5957 1716 6128 1763
rect 6540 1869 6711 1916
rect 6540 1835 6546 1869
rect 6580 1835 6711 1869
rect 6540 1797 6711 1835
rect 6540 1763 6546 1797
rect 6580 1763 6711 1797
rect 6540 1716 6711 1763
rect 5957 1416 6082 1716
rect 6138 1678 6530 1684
rect 6138 1644 6173 1678
rect 6207 1644 6245 1678
rect 6279 1644 6317 1678
rect 6351 1644 6389 1678
rect 6423 1644 6461 1678
rect 6495 1644 6530 1678
rect 6138 1593 6530 1644
rect 6138 1541 6283 1593
rect 6335 1541 6347 1593
rect 6399 1541 6530 1593
rect 6138 1488 6530 1541
rect 6138 1454 6173 1488
rect 6207 1454 6245 1488
rect 6279 1454 6317 1488
rect 6351 1454 6389 1488
rect 6423 1454 6461 1488
rect 6495 1454 6530 1488
rect 6138 1448 6530 1454
rect 6586 1416 6711 1716
rect 5957 1369 6128 1416
rect 5957 1335 6088 1369
rect 6122 1335 6128 1369
rect 5957 1297 6128 1335
rect 5957 1263 6088 1297
rect 6122 1263 6128 1297
rect 5957 1216 6128 1263
rect 6540 1369 6711 1416
rect 6540 1335 6546 1369
rect 6580 1335 6711 1369
rect 6540 1297 6711 1335
rect 6540 1263 6546 1297
rect 6580 1263 6711 1297
rect 6540 1216 6711 1263
rect 5957 1010 6082 1216
rect 6138 1178 6530 1184
rect 6138 1144 6173 1178
rect 6207 1144 6245 1178
rect 6279 1144 6317 1178
rect 6351 1144 6389 1178
rect 6423 1144 6461 1178
rect 6495 1144 6530 1178
rect 6138 1138 6530 1144
rect 5957 1009 6401 1010
rect 5957 997 6402 1009
rect 5957 963 6284 997
rect 6318 963 6356 997
rect 6390 963 6402 997
rect 5957 951 6402 963
rect 5957 943 6401 951
rect 5957 713 6082 943
rect 6586 860 6711 1216
rect 6957 2134 7403 2142
rect 6957 2100 7285 2134
rect 7319 2100 7357 2134
rect 7391 2100 7403 2134
rect 6957 2088 7403 2100
rect 6957 2075 7401 2088
rect 6957 1916 7082 2075
rect 7138 1988 7530 1994
rect 7138 1954 7173 1988
rect 7207 1954 7245 1988
rect 7279 1954 7317 1988
rect 7351 1954 7389 1988
rect 7423 1954 7461 1988
rect 7495 1954 7530 1988
rect 7138 1948 7530 1954
rect 7586 1916 7711 2397
rect 8273 2142 8403 2146
rect 6957 1869 7128 1916
rect 6957 1835 7088 1869
rect 7122 1835 7128 1869
rect 6957 1797 7128 1835
rect 6957 1763 7088 1797
rect 7122 1763 7128 1797
rect 6957 1716 7128 1763
rect 7540 1869 7711 1916
rect 7540 1835 7546 1869
rect 7580 1835 7711 1869
rect 7540 1797 7711 1835
rect 7540 1763 7546 1797
rect 7580 1763 7711 1797
rect 7540 1716 7711 1763
rect 6957 1416 7082 1716
rect 7138 1678 7530 1684
rect 7138 1644 7173 1678
rect 7207 1644 7245 1678
rect 7279 1644 7317 1678
rect 7351 1644 7389 1678
rect 7423 1644 7461 1678
rect 7495 1644 7530 1678
rect 7138 1593 7530 1644
rect 7138 1541 7283 1593
rect 7335 1541 7347 1593
rect 7399 1541 7530 1593
rect 7138 1488 7530 1541
rect 7138 1454 7173 1488
rect 7207 1454 7245 1488
rect 7279 1454 7317 1488
rect 7351 1454 7389 1488
rect 7423 1454 7461 1488
rect 7495 1454 7530 1488
rect 7138 1448 7530 1454
rect 7586 1416 7711 1716
rect 6957 1369 7128 1416
rect 6957 1335 7088 1369
rect 7122 1335 7128 1369
rect 6957 1297 7128 1335
rect 6957 1263 7088 1297
rect 7122 1263 7128 1297
rect 6957 1216 7128 1263
rect 7540 1369 7711 1416
rect 7540 1335 7546 1369
rect 7580 1335 7711 1369
rect 7540 1297 7711 1335
rect 7540 1263 7546 1297
rect 7580 1263 7711 1297
rect 7540 1216 7711 1263
rect 6957 1010 7082 1216
rect 7138 1178 7530 1184
rect 7138 1144 7173 1178
rect 7207 1144 7245 1178
rect 7279 1144 7317 1178
rect 7351 1144 7389 1178
rect 7423 1144 7461 1178
rect 7495 1144 7530 1178
rect 7138 1138 7530 1144
rect 6957 1009 7401 1010
rect 6957 997 7402 1009
rect 6957 963 7284 997
rect 7318 963 7356 997
rect 7390 963 7402 997
rect 6957 951 7402 963
rect 6957 943 7401 951
rect 6957 713 7082 943
rect 7586 860 7711 1216
rect 7957 2134 8403 2142
rect 7957 2100 8285 2134
rect 8319 2100 8357 2134
rect 8391 2100 8403 2134
rect 7957 2088 8403 2100
rect 7957 2075 8401 2088
rect 7957 1916 8082 2075
rect 8138 1988 8530 1994
rect 8138 1954 8173 1988
rect 8207 1954 8245 1988
rect 8279 1954 8317 1988
rect 8351 1954 8389 1988
rect 8423 1954 8461 1988
rect 8495 1954 8530 1988
rect 8138 1948 8530 1954
rect 8586 1916 8711 2397
rect 9273 2142 9403 2146
rect 7957 1869 8128 1916
rect 7957 1835 8088 1869
rect 8122 1835 8128 1869
rect 7957 1797 8128 1835
rect 7957 1763 8088 1797
rect 8122 1763 8128 1797
rect 7957 1716 8128 1763
rect 8540 1869 8711 1916
rect 8540 1835 8546 1869
rect 8580 1835 8711 1869
rect 8540 1797 8711 1835
rect 8540 1763 8546 1797
rect 8580 1763 8711 1797
rect 8540 1716 8711 1763
rect 7957 1416 8082 1716
rect 8138 1678 8530 1684
rect 8138 1644 8173 1678
rect 8207 1644 8245 1678
rect 8279 1644 8317 1678
rect 8351 1644 8389 1678
rect 8423 1644 8461 1678
rect 8495 1644 8530 1678
rect 8138 1593 8530 1644
rect 8138 1541 8283 1593
rect 8335 1541 8347 1593
rect 8399 1541 8530 1593
rect 8138 1488 8530 1541
rect 8138 1454 8173 1488
rect 8207 1454 8245 1488
rect 8279 1454 8317 1488
rect 8351 1454 8389 1488
rect 8423 1454 8461 1488
rect 8495 1454 8530 1488
rect 8138 1448 8530 1454
rect 8586 1416 8711 1716
rect 7957 1369 8128 1416
rect 7957 1335 8088 1369
rect 8122 1335 8128 1369
rect 7957 1297 8128 1335
rect 7957 1263 8088 1297
rect 8122 1263 8128 1297
rect 7957 1216 8128 1263
rect 8540 1369 8711 1416
rect 8540 1335 8546 1369
rect 8580 1335 8711 1369
rect 8540 1297 8711 1335
rect 8540 1263 8546 1297
rect 8580 1263 8711 1297
rect 8540 1216 8711 1263
rect 7957 1010 8082 1216
rect 8138 1178 8530 1184
rect 8138 1144 8173 1178
rect 8207 1144 8245 1178
rect 8279 1144 8317 1178
rect 8351 1144 8389 1178
rect 8423 1144 8461 1178
rect 8495 1144 8530 1178
rect 8138 1138 8530 1144
rect 7957 1009 8401 1010
rect 7957 997 8402 1009
rect 7957 963 8284 997
rect 8318 963 8356 997
rect 8390 963 8402 997
rect 7957 951 8402 963
rect 7957 943 8401 951
rect 7957 713 8082 943
rect 8586 860 8711 1216
rect 8957 2134 9403 2142
rect 8957 2100 9285 2134
rect 9319 2100 9357 2134
rect 9391 2100 9403 2134
rect 8957 2088 9403 2100
rect 8957 2075 9401 2088
rect 8957 1916 9082 2075
rect 9138 1988 9530 1994
rect 9138 1954 9173 1988
rect 9207 1954 9245 1988
rect 9279 1954 9317 1988
rect 9351 1954 9389 1988
rect 9423 1954 9461 1988
rect 9495 1954 9530 1988
rect 9138 1948 9530 1954
rect 9586 1916 9711 2397
rect 10273 2142 10403 2146
rect 8957 1869 9128 1916
rect 8957 1835 9088 1869
rect 9122 1835 9128 1869
rect 8957 1797 9128 1835
rect 8957 1763 9088 1797
rect 9122 1763 9128 1797
rect 8957 1716 9128 1763
rect 9540 1869 9711 1916
rect 9540 1835 9546 1869
rect 9580 1835 9711 1869
rect 9540 1797 9711 1835
rect 9540 1763 9546 1797
rect 9580 1763 9711 1797
rect 9540 1716 9711 1763
rect 8957 1416 9082 1716
rect 9138 1678 9530 1684
rect 9138 1644 9173 1678
rect 9207 1644 9245 1678
rect 9279 1644 9317 1678
rect 9351 1644 9389 1678
rect 9423 1644 9461 1678
rect 9495 1644 9530 1678
rect 9138 1593 9530 1644
rect 9138 1541 9283 1593
rect 9335 1541 9347 1593
rect 9399 1541 9530 1593
rect 9138 1488 9530 1541
rect 9138 1454 9173 1488
rect 9207 1454 9245 1488
rect 9279 1454 9317 1488
rect 9351 1454 9389 1488
rect 9423 1454 9461 1488
rect 9495 1454 9530 1488
rect 9138 1448 9530 1454
rect 9586 1416 9711 1716
rect 8957 1369 9128 1416
rect 8957 1335 9088 1369
rect 9122 1335 9128 1369
rect 8957 1297 9128 1335
rect 8957 1263 9088 1297
rect 9122 1263 9128 1297
rect 8957 1216 9128 1263
rect 9540 1369 9711 1416
rect 9540 1335 9546 1369
rect 9580 1335 9711 1369
rect 9540 1297 9711 1335
rect 9540 1263 9546 1297
rect 9580 1263 9711 1297
rect 9540 1216 9711 1263
rect 8957 1010 9082 1216
rect 9138 1178 9530 1184
rect 9138 1144 9173 1178
rect 9207 1144 9245 1178
rect 9279 1144 9317 1178
rect 9351 1144 9389 1178
rect 9423 1144 9461 1178
rect 9495 1144 9530 1178
rect 9138 1138 9530 1144
rect 8957 1009 9401 1010
rect 8957 997 9402 1009
rect 8957 963 9284 997
rect 9318 963 9356 997
rect 9390 963 9402 997
rect 8957 951 9402 963
rect 8957 943 9401 951
rect 8957 713 9082 943
rect 9586 860 9711 1216
rect 9957 2134 10403 2142
rect 9957 2100 10285 2134
rect 10319 2100 10357 2134
rect 10391 2100 10403 2134
rect 9957 2088 10403 2100
rect 9957 2075 10401 2088
rect 9957 1916 10082 2075
rect 10138 1988 10530 1994
rect 10138 1954 10173 1988
rect 10207 1954 10245 1988
rect 10279 1954 10317 1988
rect 10351 1954 10389 1988
rect 10423 1954 10461 1988
rect 10495 1954 10530 1988
rect 10138 1948 10530 1954
rect 10586 1916 10711 2397
rect 9957 1869 10128 1916
rect 9957 1835 10088 1869
rect 10122 1835 10128 1869
rect 9957 1797 10128 1835
rect 9957 1763 10088 1797
rect 10122 1763 10128 1797
rect 9957 1716 10128 1763
rect 10540 1869 10711 1916
rect 10540 1835 10546 1869
rect 10580 1835 10711 1869
rect 10540 1797 10711 1835
rect 10540 1763 10546 1797
rect 10580 1763 10711 1797
rect 10540 1716 10711 1763
rect 9957 1416 10082 1716
rect 10138 1678 10530 1684
rect 10138 1644 10173 1678
rect 10207 1644 10245 1678
rect 10279 1644 10317 1678
rect 10351 1644 10389 1678
rect 10423 1644 10461 1678
rect 10495 1644 10530 1678
rect 10138 1593 10530 1644
rect 10138 1541 10283 1593
rect 10335 1541 10347 1593
rect 10399 1541 10530 1593
rect 10138 1488 10530 1541
rect 10138 1454 10173 1488
rect 10207 1454 10245 1488
rect 10279 1454 10317 1488
rect 10351 1454 10389 1488
rect 10423 1454 10461 1488
rect 10495 1454 10530 1488
rect 10138 1448 10530 1454
rect 10586 1416 10711 1716
rect 9957 1369 10128 1416
rect 9957 1335 10088 1369
rect 10122 1335 10128 1369
rect 9957 1297 10128 1335
rect 9957 1263 10088 1297
rect 10122 1263 10128 1297
rect 9957 1216 10128 1263
rect 10540 1369 10711 1416
rect 10540 1335 10546 1369
rect 10580 1335 10711 1369
rect 10540 1297 10711 1335
rect 10540 1263 10546 1297
rect 10580 1263 10711 1297
rect 10540 1216 10711 1263
rect 9957 1010 10082 1216
rect 10138 1178 10530 1184
rect 10138 1144 10173 1178
rect 10207 1144 10245 1178
rect 10279 1144 10317 1178
rect 10351 1144 10389 1178
rect 10423 1144 10461 1178
rect 10495 1144 10530 1178
rect 10138 1138 10530 1144
rect 9957 1009 10401 1010
rect 9957 997 10402 1009
rect 9957 963 10284 997
rect 10318 963 10356 997
rect 10390 963 10402 997
rect 9957 951 10402 963
rect 9957 943 10401 951
rect 9957 713 10082 943
rect 10586 860 10711 1216
rect -9200 664 10818 713
rect -9200 612 -4767 664
rect -4715 612 10818 664
rect -9200 600 10818 612
rect -9200 548 -4767 600
rect -4715 548 10818 600
rect -9200 495 10818 548
rect -9200 490 -8990 495
<< via1 >>
rect 2176 7917 2228 7969
rect 2240 7917 2292 7969
rect 3176 7917 3228 7969
rect 3240 7917 3292 7969
rect 21481 8835 21533 8887
rect 21481 8771 21533 8823
rect 9938 6252 9990 6304
rect 10002 6252 10054 6304
rect -4768 5890 -4716 5942
rect -4768 5826 -4716 5878
rect 11894 6253 11946 6305
rect 11958 6253 12010 6305
rect 12794 6253 12846 6305
rect 12858 6253 12910 6305
rect 13694 6253 13746 6305
rect 13758 6253 13810 6305
rect 14594 6253 14646 6305
rect 14658 6253 14710 6305
rect 15494 6253 15546 6305
rect 15558 6253 15610 6305
rect 16394 6253 16446 6305
rect 16458 6253 16510 6305
rect 17294 6253 17346 6305
rect 17358 6253 17410 6305
rect 18194 6253 18246 6305
rect 18258 6253 18310 6305
rect 21089 5930 21141 5982
rect 21089 5866 21141 5918
rect -4165 3431 -4113 3483
rect -4101 3431 -4049 3483
rect -3465 3431 -3413 3483
rect -3401 3431 -3349 3483
rect -2765 3431 -2713 3483
rect -2701 3431 -2649 3483
rect -2065 3431 -2013 3483
rect -2001 3431 -1949 3483
rect -1365 3431 -1313 3483
rect -1301 3431 -1249 3483
rect -665 3431 -613 3483
rect -601 3431 -549 3483
rect 35 3431 87 3483
rect 99 3431 151 3483
rect 735 3431 787 3483
rect 799 3431 851 3483
rect 1435 3431 1487 3483
rect 1499 3431 1551 3483
rect 2135 3431 2187 3483
rect 2199 3431 2251 3483
rect 3835 3431 3887 3483
rect 3899 3431 3951 3483
rect 4535 3431 4587 3483
rect 4599 3431 4651 3483
rect 5235 3431 5287 3483
rect 5299 3431 5351 3483
rect 5935 3431 5987 3483
rect 5999 3431 6051 3483
rect 6635 3431 6687 3483
rect 6699 3431 6751 3483
rect 7335 3431 7387 3483
rect 7399 3431 7451 3483
rect 8035 3431 8087 3483
rect 8099 3431 8151 3483
rect 8735 3431 8787 3483
rect 8799 3431 8851 3483
rect 9435 3431 9487 3483
rect 9499 3431 9551 3483
rect 10135 3431 10187 3483
rect 10199 3431 10251 3483
rect -4767 2699 -4715 2751
rect -4767 2635 -4715 2687
rect 1283 1541 1335 1593
rect 1347 1541 1399 1593
rect 2283 1541 2335 1593
rect 2347 1541 2399 1593
rect 3283 1541 3335 1593
rect 3347 1541 3399 1593
rect 4283 1541 4335 1593
rect 4347 1541 4399 1593
rect 5283 1541 5335 1593
rect 5347 1541 5399 1593
rect 6283 1541 6335 1593
rect 6347 1541 6399 1593
rect 7283 1541 7335 1593
rect 7347 1541 7399 1593
rect 8283 1541 8335 1593
rect 8347 1541 8399 1593
rect 9283 1541 9335 1593
rect 9347 1541 9399 1593
rect 10283 1541 10335 1593
rect 10347 1541 10399 1593
rect -4767 612 -4715 664
rect -4767 548 -4715 600
<< metal2 >>
rect 11673 17085 11838 17121
rect 11673 17029 11726 17085
rect 11782 17029 11838 17085
rect 11673 17005 11838 17029
rect 11673 16949 11726 17005
rect 11782 16949 11838 17005
rect 2163 7969 3303 7979
rect 2163 7917 2176 7969
rect 2228 7917 2240 7969
rect 2292 7917 3176 7969
rect 3228 7917 3240 7969
rect 3292 7917 3303 7969
rect 2163 7904 3303 7917
rect 11673 6329 11838 16949
rect 21460 8895 21556 8905
rect 21460 8839 21478 8895
rect 21534 8839 21556 8895
rect 21460 8835 21481 8839
rect 21533 8835 21556 8839
rect 21460 8823 21556 8835
rect 21460 8815 21481 8823
rect 21533 8815 21556 8823
rect 21460 8759 21478 8815
rect 21534 8759 21556 8815
rect 21460 8743 21556 8759
rect 9880 6305 18331 6329
rect 9880 6304 11894 6305
rect 9880 6252 9938 6304
rect 9990 6252 10002 6304
rect 10054 6253 11894 6304
rect 11946 6253 11958 6305
rect 12010 6253 12794 6305
rect 12846 6253 12858 6305
rect 12910 6253 13694 6305
rect 13746 6253 13758 6305
rect 13810 6253 14594 6305
rect 14646 6253 14658 6305
rect 14710 6253 15494 6305
rect 15546 6253 15558 6305
rect 15610 6253 16394 6305
rect 16446 6253 16458 6305
rect 16510 6253 17294 6305
rect 17346 6253 17358 6305
rect 17410 6253 18194 6305
rect 18246 6253 18258 6305
rect 18310 6253 18331 6305
rect 10054 6252 18331 6253
rect 9880 6229 18331 6252
rect 21083 5982 21147 5988
rect 21083 5953 21089 5982
rect -4794 5942 21089 5953
rect -4794 5890 -4768 5942
rect -4716 5930 21089 5942
rect 21141 5953 21147 5982
rect 21141 5930 21155 5953
rect -4716 5918 21155 5930
rect -4716 5890 21089 5918
rect -4794 5878 21089 5890
rect -4794 5853 -4768 5878
rect -4774 5826 -4768 5853
rect -4716 5866 21089 5878
rect 21141 5866 21155 5918
rect -4716 5853 21155 5866
rect -4716 5826 -4710 5853
rect -4774 5820 -4710 5826
rect -9200 3499 -9040 3500
rect -9200 3483 2273 3499
rect -9200 3431 -4165 3483
rect -4113 3431 -4101 3483
rect -4049 3431 -3465 3483
rect -3413 3431 -3401 3483
rect -3349 3431 -2765 3483
rect -2713 3431 -2701 3483
rect -2649 3431 -2065 3483
rect -2013 3431 -2001 3483
rect -1949 3431 -1365 3483
rect -1313 3431 -1301 3483
rect -1249 3431 -665 3483
rect -613 3431 -601 3483
rect -549 3431 35 3483
rect 87 3431 99 3483
rect 151 3431 735 3483
rect 787 3431 799 3483
rect 851 3431 1435 3483
rect 1487 3431 1499 3483
rect 1551 3431 2135 3483
rect 2187 3431 2199 3483
rect 2251 3431 2273 3483
rect -9200 3414 2273 3431
rect 3819 3483 33850 3499
rect 3819 3431 3835 3483
rect 3887 3431 3899 3483
rect 3951 3431 4535 3483
rect 4587 3431 4599 3483
rect 4651 3431 5235 3483
rect 5287 3431 5299 3483
rect 5351 3431 5935 3483
rect 5987 3431 5999 3483
rect 6051 3431 6635 3483
rect 6687 3431 6699 3483
rect 6751 3431 7335 3483
rect 7387 3431 7399 3483
rect 7451 3431 8035 3483
rect 8087 3431 8099 3483
rect 8151 3431 8735 3483
rect 8787 3431 8799 3483
rect 8851 3431 9435 3483
rect 9487 3431 9499 3483
rect 9551 3431 10135 3483
rect 10187 3431 10199 3483
rect 10251 3431 33850 3483
rect 3819 3414 33850 3431
rect -9200 3410 -9040 3414
rect -4780 2751 -4702 2762
rect -4780 2699 -4767 2751
rect -4715 2699 -4702 2751
rect -4780 2687 -4702 2699
rect -4780 2635 -4767 2687
rect -4715 2635 -4702 2687
rect -4780 664 -4702 2635
rect 1268 1593 10427 1609
rect 1268 1541 1283 1593
rect 1335 1541 1347 1593
rect 1399 1541 2283 1593
rect 2335 1541 2347 1593
rect 2399 1541 3283 1593
rect 3335 1541 3347 1593
rect 3399 1541 4283 1593
rect 4335 1541 4347 1593
rect 4399 1541 5283 1593
rect 5335 1541 5347 1593
rect 5399 1541 6283 1593
rect 6335 1541 6347 1593
rect 6399 1541 7283 1593
rect 7335 1541 7347 1593
rect 7399 1541 8283 1593
rect 8335 1541 8347 1593
rect 8399 1541 9283 1593
rect 9335 1541 9347 1593
rect 9399 1541 10283 1593
rect 10335 1541 10347 1593
rect 10399 1541 10427 1593
rect 1268 1525 10427 1541
rect -4780 612 -4767 664
rect -4715 612 -4702 664
rect -4780 600 -4702 612
rect -4780 548 -4767 600
rect -4715 548 -4702 600
rect -4780 507 -4702 548
<< via2 >>
rect 11726 17029 11782 17085
rect 11726 16949 11782 17005
rect 21478 8887 21534 8895
rect 21478 8839 21481 8887
rect 21481 8839 21533 8887
rect 21533 8839 21534 8887
rect 21478 8771 21481 8815
rect 21481 8771 21533 8815
rect 21533 8771 21534 8815
rect 21478 8759 21534 8771
<< metal3 >>
rect 11718 17107 11794 17112
rect 11707 17106 11804 17107
rect 11707 17042 11724 17106
rect 11788 17042 11804 17106
rect 11707 17029 11726 17042
rect 11782 17029 11804 17042
rect 11707 17005 11804 17029
rect 11707 16996 11726 17005
rect 11782 16996 11804 17005
rect 11707 16932 11724 16996
rect 11788 16932 11804 16996
rect 11707 16925 11804 16932
rect -8719 10453 -2519 16668
rect -8719 10389 -8691 10453
rect -8627 10389 -8611 10453
rect -8547 10389 -8531 10453
rect -8467 10389 -8451 10453
rect -8387 10389 -8371 10453
rect -8307 10389 -8291 10453
rect -8227 10389 -8211 10453
rect -8147 10389 -8131 10453
rect -8067 10389 -8051 10453
rect -7987 10389 -7971 10453
rect -7907 10389 -7891 10453
rect -7827 10389 -7811 10453
rect -7747 10389 -7731 10453
rect -7667 10389 -7651 10453
rect -7587 10389 -7571 10453
rect -7507 10389 -7491 10453
rect -7427 10389 -7411 10453
rect -7347 10389 -7331 10453
rect -7267 10389 -7251 10453
rect -7187 10389 -7171 10453
rect -7107 10389 -7091 10453
rect -7027 10389 -7011 10453
rect -6947 10389 -6931 10453
rect -6867 10389 -6851 10453
rect -6787 10389 -6771 10453
rect -6707 10389 -6691 10453
rect -6627 10389 -6611 10453
rect -6547 10389 -6531 10453
rect -6467 10389 -6451 10453
rect -6387 10389 -6371 10453
rect -6307 10389 -6291 10453
rect -6227 10389 -6211 10453
rect -6147 10389 -6131 10453
rect -6067 10389 -6051 10453
rect -5987 10389 -5971 10453
rect -5907 10389 -5891 10453
rect -5827 10389 -5811 10453
rect -5747 10389 -5731 10453
rect -5667 10389 -5651 10453
rect -5587 10389 -5571 10453
rect -5507 10389 -5491 10453
rect -5427 10389 -5411 10453
rect -5347 10389 -5331 10453
rect -5267 10389 -5251 10453
rect -5187 10389 -5171 10453
rect -5107 10389 -5091 10453
rect -5027 10389 -5011 10453
rect -4947 10389 -4931 10453
rect -4867 10389 -4851 10453
rect -4787 10389 -4771 10453
rect -4707 10389 -4691 10453
rect -4627 10389 -4611 10453
rect -4547 10389 -4531 10453
rect -4467 10389 -4451 10453
rect -4387 10389 -4371 10453
rect -4307 10389 -4291 10453
rect -4227 10389 -4211 10453
rect -4147 10389 -4131 10453
rect -4067 10389 -4051 10453
rect -3987 10389 -3971 10453
rect -3907 10389 -3891 10453
rect -3827 10389 -3811 10453
rect -3747 10389 -3731 10453
rect -3667 10389 -3651 10453
rect -3587 10389 -3571 10453
rect -3507 10389 -3491 10453
rect -3427 10389 -3411 10453
rect -3347 10389 -3331 10453
rect -3267 10389 -3251 10453
rect -3187 10389 -3171 10453
rect -3107 10389 -3091 10453
rect -3027 10389 -3011 10453
rect -2947 10389 -2931 10453
rect -2867 10389 -2851 10453
rect -2787 10389 -2771 10453
rect -2707 10389 -2691 10453
rect -2627 10389 -2611 10453
rect -2547 10389 -2519 10453
rect -8719 10369 -2519 10389
rect -1719 10453 4481 16668
rect -1719 10389 -1691 10453
rect -1627 10389 -1611 10453
rect -1547 10389 -1531 10453
rect -1467 10389 -1451 10453
rect -1387 10389 -1371 10453
rect -1307 10389 -1291 10453
rect -1227 10389 -1211 10453
rect -1147 10389 -1131 10453
rect -1067 10389 -1051 10453
rect -987 10389 -971 10453
rect -907 10389 -891 10453
rect -827 10389 -811 10453
rect -747 10389 -731 10453
rect -667 10389 -651 10453
rect -587 10389 -571 10453
rect -507 10389 -491 10453
rect -427 10389 -411 10453
rect -347 10389 -331 10453
rect -267 10389 -251 10453
rect -187 10389 -171 10453
rect -107 10389 -91 10453
rect -27 10389 -11 10453
rect 53 10389 69 10453
rect 133 10389 149 10453
rect 213 10389 229 10453
rect 293 10389 309 10453
rect 373 10389 389 10453
rect 453 10389 469 10453
rect 533 10389 549 10453
rect 613 10389 629 10453
rect 693 10389 709 10453
rect 773 10389 789 10453
rect 853 10389 869 10453
rect 933 10389 949 10453
rect 1013 10389 1029 10453
rect 1093 10389 1109 10453
rect 1173 10389 1189 10453
rect 1253 10389 1269 10453
rect 1333 10389 1349 10453
rect 1413 10389 1429 10453
rect 1493 10389 1509 10453
rect 1573 10389 1589 10453
rect 1653 10389 1669 10453
rect 1733 10389 1749 10453
rect 1813 10389 1829 10453
rect 1893 10389 1909 10453
rect 1973 10389 1989 10453
rect 2053 10389 2069 10453
rect 2133 10389 2149 10453
rect 2213 10389 2229 10453
rect 2293 10389 2309 10453
rect 2373 10389 2389 10453
rect 2453 10389 2469 10453
rect 2533 10389 2549 10453
rect 2613 10389 2629 10453
rect 2693 10389 2709 10453
rect 2773 10389 2789 10453
rect 2853 10389 2869 10453
rect 2933 10389 2949 10453
rect 3013 10389 3029 10453
rect 3093 10389 3109 10453
rect 3173 10389 3189 10453
rect 3253 10389 3269 10453
rect 3333 10389 3349 10453
rect 3413 10389 3429 10453
rect 3493 10389 3509 10453
rect 3573 10389 3589 10453
rect 3653 10389 3669 10453
rect 3733 10389 3749 10453
rect 3813 10389 3829 10453
rect 3893 10389 3909 10453
rect 3973 10389 3989 10453
rect 4053 10389 4069 10453
rect 4133 10389 4149 10453
rect 4213 10389 4229 10453
rect 4293 10389 4309 10453
rect 4373 10389 4389 10453
rect 4453 10389 4481 10453
rect -1719 10369 4481 10389
rect 5281 10453 11481 16668
rect 5281 10389 5309 10453
rect 5373 10389 5389 10453
rect 5453 10389 5469 10453
rect 5533 10389 5549 10453
rect 5613 10389 5629 10453
rect 5693 10389 5709 10453
rect 5773 10389 5789 10453
rect 5853 10389 5869 10453
rect 5933 10389 5949 10453
rect 6013 10389 6029 10453
rect 6093 10389 6109 10453
rect 6173 10389 6189 10453
rect 6253 10389 6269 10453
rect 6333 10389 6349 10453
rect 6413 10389 6429 10453
rect 6493 10389 6509 10453
rect 6573 10389 6589 10453
rect 6653 10389 6669 10453
rect 6733 10389 6749 10453
rect 6813 10389 6829 10453
rect 6893 10389 6909 10453
rect 6973 10389 6989 10453
rect 7053 10389 7069 10453
rect 7133 10389 7149 10453
rect 7213 10389 7229 10453
rect 7293 10389 7309 10453
rect 7373 10389 7389 10453
rect 7453 10389 7469 10453
rect 7533 10389 7549 10453
rect 7613 10389 7629 10453
rect 7693 10389 7709 10453
rect 7773 10389 7789 10453
rect 7853 10389 7869 10453
rect 7933 10389 7949 10453
rect 8013 10389 8029 10453
rect 8093 10389 8109 10453
rect 8173 10389 8189 10453
rect 8253 10389 8269 10453
rect 8333 10389 8349 10453
rect 8413 10389 8429 10453
rect 8493 10389 8509 10453
rect 8573 10389 8589 10453
rect 8653 10389 8669 10453
rect 8733 10389 8749 10453
rect 8813 10389 8829 10453
rect 8893 10389 8909 10453
rect 8973 10389 8989 10453
rect 9053 10389 9069 10453
rect 9133 10389 9149 10453
rect 9213 10389 9229 10453
rect 9293 10389 9309 10453
rect 9373 10389 9389 10453
rect 9453 10389 9469 10453
rect 9533 10389 9549 10453
rect 9613 10389 9629 10453
rect 9693 10389 9709 10453
rect 9773 10389 9789 10453
rect 9853 10389 9869 10453
rect 9933 10389 9949 10453
rect 10013 10389 10029 10453
rect 10093 10389 10109 10453
rect 10173 10389 10189 10453
rect 10253 10389 10269 10453
rect 10333 10389 10349 10453
rect 10413 10389 10429 10453
rect 10493 10389 10509 10453
rect 10573 10389 10589 10453
rect 10653 10389 10669 10453
rect 10733 10389 10749 10453
rect 10813 10389 10829 10453
rect 10893 10389 10909 10453
rect 10973 10389 10989 10453
rect 11053 10389 11069 10453
rect 11133 10389 11149 10453
rect 11213 10389 11229 10453
rect 11293 10389 11309 10453
rect 11373 10389 11389 10453
rect 11453 10389 11481 10453
rect 5281 10369 11481 10389
rect 12281 10453 18481 16668
rect 12281 10389 12309 10453
rect 12373 10389 12389 10453
rect 12453 10389 12469 10453
rect 12533 10389 12549 10453
rect 12613 10389 12629 10453
rect 12693 10389 12709 10453
rect 12773 10389 12789 10453
rect 12853 10389 12869 10453
rect 12933 10389 12949 10453
rect 13013 10389 13029 10453
rect 13093 10389 13109 10453
rect 13173 10389 13189 10453
rect 13253 10389 13269 10453
rect 13333 10389 13349 10453
rect 13413 10389 13429 10453
rect 13493 10389 13509 10453
rect 13573 10389 13589 10453
rect 13653 10389 13669 10453
rect 13733 10389 13749 10453
rect 13813 10389 13829 10453
rect 13893 10389 13909 10453
rect 13973 10389 13989 10453
rect 14053 10389 14069 10453
rect 14133 10389 14149 10453
rect 14213 10389 14229 10453
rect 14293 10389 14309 10453
rect 14373 10389 14389 10453
rect 14453 10389 14469 10453
rect 14533 10389 14549 10453
rect 14613 10389 14629 10453
rect 14693 10389 14709 10453
rect 14773 10389 14789 10453
rect 14853 10389 14869 10453
rect 14933 10389 14949 10453
rect 15013 10389 15029 10453
rect 15093 10389 15109 10453
rect 15173 10389 15189 10453
rect 15253 10389 15269 10453
rect 15333 10389 15349 10453
rect 15413 10389 15429 10453
rect 15493 10389 15509 10453
rect 15573 10389 15589 10453
rect 15653 10389 15669 10453
rect 15733 10389 15749 10453
rect 15813 10389 15829 10453
rect 15893 10389 15909 10453
rect 15973 10389 15989 10453
rect 16053 10389 16069 10453
rect 16133 10389 16149 10453
rect 16213 10389 16229 10453
rect 16293 10389 16309 10453
rect 16373 10389 16389 10453
rect 16453 10389 16469 10453
rect 16533 10389 16549 10453
rect 16613 10389 16629 10453
rect 16693 10389 16709 10453
rect 16773 10389 16789 10453
rect 16853 10389 16869 10453
rect 16933 10389 16949 10453
rect 17013 10389 17029 10453
rect 17093 10389 17109 10453
rect 17173 10389 17189 10453
rect 17253 10389 17269 10453
rect 17333 10389 17349 10453
rect 17413 10389 17429 10453
rect 17493 10389 17509 10453
rect 17573 10389 17589 10453
rect 17653 10389 17669 10453
rect 17733 10389 17749 10453
rect 17813 10389 17829 10453
rect 17893 10389 17909 10453
rect 17973 10389 17989 10453
rect 18053 10389 18069 10453
rect 18133 10389 18149 10453
rect 18213 10389 18229 10453
rect 18293 10389 18309 10453
rect 18373 10389 18389 10453
rect 18453 10389 18481 10453
rect 12281 10369 18481 10389
rect 19281 10453 25481 16668
rect 19281 10389 19309 10453
rect 19373 10389 19389 10453
rect 19453 10389 19469 10453
rect 19533 10389 19549 10453
rect 19613 10389 19629 10453
rect 19693 10389 19709 10453
rect 19773 10389 19789 10453
rect 19853 10389 19869 10453
rect 19933 10389 19949 10453
rect 20013 10389 20029 10453
rect 20093 10389 20109 10453
rect 20173 10389 20189 10453
rect 20253 10389 20269 10453
rect 20333 10389 20349 10453
rect 20413 10389 20429 10453
rect 20493 10389 20509 10453
rect 20573 10389 20589 10453
rect 20653 10389 20669 10453
rect 20733 10389 20749 10453
rect 20813 10389 20829 10453
rect 20893 10389 20909 10453
rect 20973 10389 20989 10453
rect 21053 10389 21069 10453
rect 21133 10389 21149 10453
rect 21213 10389 21229 10453
rect 21293 10389 21309 10453
rect 21373 10389 21389 10453
rect 21453 10389 21469 10453
rect 21533 10389 21549 10453
rect 21613 10389 21629 10453
rect 21693 10389 21709 10453
rect 21773 10389 21789 10453
rect 21853 10389 21869 10453
rect 21933 10389 21949 10453
rect 22013 10389 22029 10453
rect 22093 10389 22109 10453
rect 22173 10389 22189 10453
rect 22253 10389 22269 10453
rect 22333 10389 22349 10453
rect 22413 10389 22429 10453
rect 22493 10389 22509 10453
rect 22573 10389 22589 10453
rect 22653 10389 22669 10453
rect 22733 10389 22749 10453
rect 22813 10389 22829 10453
rect 22893 10389 22909 10453
rect 22973 10389 22989 10453
rect 23053 10389 23069 10453
rect 23133 10389 23149 10453
rect 23213 10389 23229 10453
rect 23293 10389 23309 10453
rect 23373 10389 23389 10453
rect 23453 10389 23469 10453
rect 23533 10389 23549 10453
rect 23613 10389 23629 10453
rect 23693 10389 23709 10453
rect 23773 10389 23789 10453
rect 23853 10389 23869 10453
rect 23933 10389 23949 10453
rect 24013 10389 24029 10453
rect 24093 10389 24109 10453
rect 24173 10389 24189 10453
rect 24253 10389 24269 10453
rect 24333 10389 24349 10453
rect 24413 10389 24429 10453
rect 24493 10389 24509 10453
rect 24573 10389 24589 10453
rect 24653 10389 24669 10453
rect 24733 10389 24749 10453
rect 24813 10389 24829 10453
rect 24893 10389 24909 10453
rect 24973 10389 24989 10453
rect 25053 10389 25069 10453
rect 25133 10389 25149 10453
rect 25213 10389 25229 10453
rect 25293 10389 25309 10453
rect 25373 10389 25389 10453
rect 25453 10389 25481 10453
rect 19281 10369 25481 10389
rect 26281 10453 32481 16668
rect 26281 10389 26309 10453
rect 26373 10389 26389 10453
rect 26453 10389 26469 10453
rect 26533 10389 26549 10453
rect 26613 10389 26629 10453
rect 26693 10389 26709 10453
rect 26773 10389 26789 10453
rect 26853 10389 26869 10453
rect 26933 10389 26949 10453
rect 27013 10389 27029 10453
rect 27093 10389 27109 10453
rect 27173 10389 27189 10453
rect 27253 10389 27269 10453
rect 27333 10389 27349 10453
rect 27413 10389 27429 10453
rect 27493 10389 27509 10453
rect 27573 10389 27589 10453
rect 27653 10389 27669 10453
rect 27733 10389 27749 10453
rect 27813 10389 27829 10453
rect 27893 10389 27909 10453
rect 27973 10389 27989 10453
rect 28053 10389 28069 10453
rect 28133 10389 28149 10453
rect 28213 10389 28229 10453
rect 28293 10389 28309 10453
rect 28373 10389 28389 10453
rect 28453 10389 28469 10453
rect 28533 10389 28549 10453
rect 28613 10389 28629 10453
rect 28693 10389 28709 10453
rect 28773 10389 28789 10453
rect 28853 10389 28869 10453
rect 28933 10389 28949 10453
rect 29013 10389 29029 10453
rect 29093 10389 29109 10453
rect 29173 10389 29189 10453
rect 29253 10389 29269 10453
rect 29333 10389 29349 10453
rect 29413 10389 29429 10453
rect 29493 10389 29509 10453
rect 29573 10389 29589 10453
rect 29653 10389 29669 10453
rect 29733 10389 29749 10453
rect 29813 10389 29829 10453
rect 29893 10389 29909 10453
rect 29973 10389 29989 10453
rect 30053 10389 30069 10453
rect 30133 10389 30149 10453
rect 30213 10389 30229 10453
rect 30293 10389 30309 10453
rect 30373 10389 30389 10453
rect 30453 10389 30469 10453
rect 30533 10389 30549 10453
rect 30613 10389 30629 10453
rect 30693 10389 30709 10453
rect 30773 10389 30789 10453
rect 30853 10389 30869 10453
rect 30933 10389 30949 10453
rect 31013 10389 31029 10453
rect 31093 10389 31109 10453
rect 31173 10389 31189 10453
rect 31253 10389 31269 10453
rect 31333 10389 31349 10453
rect 31413 10389 31429 10453
rect 31493 10389 31509 10453
rect 31573 10389 31589 10453
rect 31653 10389 31669 10453
rect 31733 10389 31749 10453
rect 31813 10389 31829 10453
rect 31893 10389 31909 10453
rect 31973 10389 31989 10453
rect 32053 10389 32069 10453
rect 32133 10389 32149 10453
rect 32213 10389 32229 10453
rect 32293 10389 32309 10453
rect 32373 10389 32389 10453
rect 32453 10389 32481 10453
rect 26281 10369 32481 10389
rect 21470 8910 21546 8916
rect 21470 8907 21476 8910
rect 21458 8846 21476 8907
rect 21540 8907 21546 8910
rect 21540 8846 21558 8907
rect 21458 8839 21478 8846
rect 21534 8839 21558 8846
rect 21458 8815 21558 8839
rect 21458 8800 21478 8815
rect 21534 8800 21558 8815
rect 21458 8740 21476 8800
rect 21470 8736 21476 8740
rect 21540 8740 21558 8800
rect 21540 8736 21546 8740
rect 21470 8730 21546 8736
<< via3 >>
rect 11724 17085 11788 17106
rect 11724 17042 11726 17085
rect 11726 17042 11782 17085
rect 11782 17042 11788 17085
rect 11724 16949 11726 16996
rect 11726 16949 11782 16996
rect 11782 16949 11788 16996
rect 11724 16932 11788 16949
rect -8691 10389 -8627 10453
rect -8611 10389 -8547 10453
rect -8531 10389 -8467 10453
rect -8451 10389 -8387 10453
rect -8371 10389 -8307 10453
rect -8291 10389 -8227 10453
rect -8211 10389 -8147 10453
rect -8131 10389 -8067 10453
rect -8051 10389 -7987 10453
rect -7971 10389 -7907 10453
rect -7891 10389 -7827 10453
rect -7811 10389 -7747 10453
rect -7731 10389 -7667 10453
rect -7651 10389 -7587 10453
rect -7571 10389 -7507 10453
rect -7491 10389 -7427 10453
rect -7411 10389 -7347 10453
rect -7331 10389 -7267 10453
rect -7251 10389 -7187 10453
rect -7171 10389 -7107 10453
rect -7091 10389 -7027 10453
rect -7011 10389 -6947 10453
rect -6931 10389 -6867 10453
rect -6851 10389 -6787 10453
rect -6771 10389 -6707 10453
rect -6691 10389 -6627 10453
rect -6611 10389 -6547 10453
rect -6531 10389 -6467 10453
rect -6451 10389 -6387 10453
rect -6371 10389 -6307 10453
rect -6291 10389 -6227 10453
rect -6211 10389 -6147 10453
rect -6131 10389 -6067 10453
rect -6051 10389 -5987 10453
rect -5971 10389 -5907 10453
rect -5891 10389 -5827 10453
rect -5811 10389 -5747 10453
rect -5731 10389 -5667 10453
rect -5651 10389 -5587 10453
rect -5571 10389 -5507 10453
rect -5491 10389 -5427 10453
rect -5411 10389 -5347 10453
rect -5331 10389 -5267 10453
rect -5251 10389 -5187 10453
rect -5171 10389 -5107 10453
rect -5091 10389 -5027 10453
rect -5011 10389 -4947 10453
rect -4931 10389 -4867 10453
rect -4851 10389 -4787 10453
rect -4771 10389 -4707 10453
rect -4691 10389 -4627 10453
rect -4611 10389 -4547 10453
rect -4531 10389 -4467 10453
rect -4451 10389 -4387 10453
rect -4371 10389 -4307 10453
rect -4291 10389 -4227 10453
rect -4211 10389 -4147 10453
rect -4131 10389 -4067 10453
rect -4051 10389 -3987 10453
rect -3971 10389 -3907 10453
rect -3891 10389 -3827 10453
rect -3811 10389 -3747 10453
rect -3731 10389 -3667 10453
rect -3651 10389 -3587 10453
rect -3571 10389 -3507 10453
rect -3491 10389 -3427 10453
rect -3411 10389 -3347 10453
rect -3331 10389 -3267 10453
rect -3251 10389 -3187 10453
rect -3171 10389 -3107 10453
rect -3091 10389 -3027 10453
rect -3011 10389 -2947 10453
rect -2931 10389 -2867 10453
rect -2851 10389 -2787 10453
rect -2771 10389 -2707 10453
rect -2691 10389 -2627 10453
rect -2611 10389 -2547 10453
rect -1691 10389 -1627 10453
rect -1611 10389 -1547 10453
rect -1531 10389 -1467 10453
rect -1451 10389 -1387 10453
rect -1371 10389 -1307 10453
rect -1291 10389 -1227 10453
rect -1211 10389 -1147 10453
rect -1131 10389 -1067 10453
rect -1051 10389 -987 10453
rect -971 10389 -907 10453
rect -891 10389 -827 10453
rect -811 10389 -747 10453
rect -731 10389 -667 10453
rect -651 10389 -587 10453
rect -571 10389 -507 10453
rect -491 10389 -427 10453
rect -411 10389 -347 10453
rect -331 10389 -267 10453
rect -251 10389 -187 10453
rect -171 10389 -107 10453
rect -91 10389 -27 10453
rect -11 10389 53 10453
rect 69 10389 133 10453
rect 149 10389 213 10453
rect 229 10389 293 10453
rect 309 10389 373 10453
rect 389 10389 453 10453
rect 469 10389 533 10453
rect 549 10389 613 10453
rect 629 10389 693 10453
rect 709 10389 773 10453
rect 789 10389 853 10453
rect 869 10389 933 10453
rect 949 10389 1013 10453
rect 1029 10389 1093 10453
rect 1109 10389 1173 10453
rect 1189 10389 1253 10453
rect 1269 10389 1333 10453
rect 1349 10389 1413 10453
rect 1429 10389 1493 10453
rect 1509 10389 1573 10453
rect 1589 10389 1653 10453
rect 1669 10389 1733 10453
rect 1749 10389 1813 10453
rect 1829 10389 1893 10453
rect 1909 10389 1973 10453
rect 1989 10389 2053 10453
rect 2069 10389 2133 10453
rect 2149 10389 2213 10453
rect 2229 10389 2293 10453
rect 2309 10389 2373 10453
rect 2389 10389 2453 10453
rect 2469 10389 2533 10453
rect 2549 10389 2613 10453
rect 2629 10389 2693 10453
rect 2709 10389 2773 10453
rect 2789 10389 2853 10453
rect 2869 10389 2933 10453
rect 2949 10389 3013 10453
rect 3029 10389 3093 10453
rect 3109 10389 3173 10453
rect 3189 10389 3253 10453
rect 3269 10389 3333 10453
rect 3349 10389 3413 10453
rect 3429 10389 3493 10453
rect 3509 10389 3573 10453
rect 3589 10389 3653 10453
rect 3669 10389 3733 10453
rect 3749 10389 3813 10453
rect 3829 10389 3893 10453
rect 3909 10389 3973 10453
rect 3989 10389 4053 10453
rect 4069 10389 4133 10453
rect 4149 10389 4213 10453
rect 4229 10389 4293 10453
rect 4309 10389 4373 10453
rect 4389 10389 4453 10453
rect 5309 10389 5373 10453
rect 5389 10389 5453 10453
rect 5469 10389 5533 10453
rect 5549 10389 5613 10453
rect 5629 10389 5693 10453
rect 5709 10389 5773 10453
rect 5789 10389 5853 10453
rect 5869 10389 5933 10453
rect 5949 10389 6013 10453
rect 6029 10389 6093 10453
rect 6109 10389 6173 10453
rect 6189 10389 6253 10453
rect 6269 10389 6333 10453
rect 6349 10389 6413 10453
rect 6429 10389 6493 10453
rect 6509 10389 6573 10453
rect 6589 10389 6653 10453
rect 6669 10389 6733 10453
rect 6749 10389 6813 10453
rect 6829 10389 6893 10453
rect 6909 10389 6973 10453
rect 6989 10389 7053 10453
rect 7069 10389 7133 10453
rect 7149 10389 7213 10453
rect 7229 10389 7293 10453
rect 7309 10389 7373 10453
rect 7389 10389 7453 10453
rect 7469 10389 7533 10453
rect 7549 10389 7613 10453
rect 7629 10389 7693 10453
rect 7709 10389 7773 10453
rect 7789 10389 7853 10453
rect 7869 10389 7933 10453
rect 7949 10389 8013 10453
rect 8029 10389 8093 10453
rect 8109 10389 8173 10453
rect 8189 10389 8253 10453
rect 8269 10389 8333 10453
rect 8349 10389 8413 10453
rect 8429 10389 8493 10453
rect 8509 10389 8573 10453
rect 8589 10389 8653 10453
rect 8669 10389 8733 10453
rect 8749 10389 8813 10453
rect 8829 10389 8893 10453
rect 8909 10389 8973 10453
rect 8989 10389 9053 10453
rect 9069 10389 9133 10453
rect 9149 10389 9213 10453
rect 9229 10389 9293 10453
rect 9309 10389 9373 10453
rect 9389 10389 9453 10453
rect 9469 10389 9533 10453
rect 9549 10389 9613 10453
rect 9629 10389 9693 10453
rect 9709 10389 9773 10453
rect 9789 10389 9853 10453
rect 9869 10389 9933 10453
rect 9949 10389 10013 10453
rect 10029 10389 10093 10453
rect 10109 10389 10173 10453
rect 10189 10389 10253 10453
rect 10269 10389 10333 10453
rect 10349 10389 10413 10453
rect 10429 10389 10493 10453
rect 10509 10389 10573 10453
rect 10589 10389 10653 10453
rect 10669 10389 10733 10453
rect 10749 10389 10813 10453
rect 10829 10389 10893 10453
rect 10909 10389 10973 10453
rect 10989 10389 11053 10453
rect 11069 10389 11133 10453
rect 11149 10389 11213 10453
rect 11229 10389 11293 10453
rect 11309 10389 11373 10453
rect 11389 10389 11453 10453
rect 12309 10389 12373 10453
rect 12389 10389 12453 10453
rect 12469 10389 12533 10453
rect 12549 10389 12613 10453
rect 12629 10389 12693 10453
rect 12709 10389 12773 10453
rect 12789 10389 12853 10453
rect 12869 10389 12933 10453
rect 12949 10389 13013 10453
rect 13029 10389 13093 10453
rect 13109 10389 13173 10453
rect 13189 10389 13253 10453
rect 13269 10389 13333 10453
rect 13349 10389 13413 10453
rect 13429 10389 13493 10453
rect 13509 10389 13573 10453
rect 13589 10389 13653 10453
rect 13669 10389 13733 10453
rect 13749 10389 13813 10453
rect 13829 10389 13893 10453
rect 13909 10389 13973 10453
rect 13989 10389 14053 10453
rect 14069 10389 14133 10453
rect 14149 10389 14213 10453
rect 14229 10389 14293 10453
rect 14309 10389 14373 10453
rect 14389 10389 14453 10453
rect 14469 10389 14533 10453
rect 14549 10389 14613 10453
rect 14629 10389 14693 10453
rect 14709 10389 14773 10453
rect 14789 10389 14853 10453
rect 14869 10389 14933 10453
rect 14949 10389 15013 10453
rect 15029 10389 15093 10453
rect 15109 10389 15173 10453
rect 15189 10389 15253 10453
rect 15269 10389 15333 10453
rect 15349 10389 15413 10453
rect 15429 10389 15493 10453
rect 15509 10389 15573 10453
rect 15589 10389 15653 10453
rect 15669 10389 15733 10453
rect 15749 10389 15813 10453
rect 15829 10389 15893 10453
rect 15909 10389 15973 10453
rect 15989 10389 16053 10453
rect 16069 10389 16133 10453
rect 16149 10389 16213 10453
rect 16229 10389 16293 10453
rect 16309 10389 16373 10453
rect 16389 10389 16453 10453
rect 16469 10389 16533 10453
rect 16549 10389 16613 10453
rect 16629 10389 16693 10453
rect 16709 10389 16773 10453
rect 16789 10389 16853 10453
rect 16869 10389 16933 10453
rect 16949 10389 17013 10453
rect 17029 10389 17093 10453
rect 17109 10389 17173 10453
rect 17189 10389 17253 10453
rect 17269 10389 17333 10453
rect 17349 10389 17413 10453
rect 17429 10389 17493 10453
rect 17509 10389 17573 10453
rect 17589 10389 17653 10453
rect 17669 10389 17733 10453
rect 17749 10389 17813 10453
rect 17829 10389 17893 10453
rect 17909 10389 17973 10453
rect 17989 10389 18053 10453
rect 18069 10389 18133 10453
rect 18149 10389 18213 10453
rect 18229 10389 18293 10453
rect 18309 10389 18373 10453
rect 18389 10389 18453 10453
rect 19309 10389 19373 10453
rect 19389 10389 19453 10453
rect 19469 10389 19533 10453
rect 19549 10389 19613 10453
rect 19629 10389 19693 10453
rect 19709 10389 19773 10453
rect 19789 10389 19853 10453
rect 19869 10389 19933 10453
rect 19949 10389 20013 10453
rect 20029 10389 20093 10453
rect 20109 10389 20173 10453
rect 20189 10389 20253 10453
rect 20269 10389 20333 10453
rect 20349 10389 20413 10453
rect 20429 10389 20493 10453
rect 20509 10389 20573 10453
rect 20589 10389 20653 10453
rect 20669 10389 20733 10453
rect 20749 10389 20813 10453
rect 20829 10389 20893 10453
rect 20909 10389 20973 10453
rect 20989 10389 21053 10453
rect 21069 10389 21133 10453
rect 21149 10389 21213 10453
rect 21229 10389 21293 10453
rect 21309 10389 21373 10453
rect 21389 10389 21453 10453
rect 21469 10389 21533 10453
rect 21549 10389 21613 10453
rect 21629 10389 21693 10453
rect 21709 10389 21773 10453
rect 21789 10389 21853 10453
rect 21869 10389 21933 10453
rect 21949 10389 22013 10453
rect 22029 10389 22093 10453
rect 22109 10389 22173 10453
rect 22189 10389 22253 10453
rect 22269 10389 22333 10453
rect 22349 10389 22413 10453
rect 22429 10389 22493 10453
rect 22509 10389 22573 10453
rect 22589 10389 22653 10453
rect 22669 10389 22733 10453
rect 22749 10389 22813 10453
rect 22829 10389 22893 10453
rect 22909 10389 22973 10453
rect 22989 10389 23053 10453
rect 23069 10389 23133 10453
rect 23149 10389 23213 10453
rect 23229 10389 23293 10453
rect 23309 10389 23373 10453
rect 23389 10389 23453 10453
rect 23469 10389 23533 10453
rect 23549 10389 23613 10453
rect 23629 10389 23693 10453
rect 23709 10389 23773 10453
rect 23789 10389 23853 10453
rect 23869 10389 23933 10453
rect 23949 10389 24013 10453
rect 24029 10389 24093 10453
rect 24109 10389 24173 10453
rect 24189 10389 24253 10453
rect 24269 10389 24333 10453
rect 24349 10389 24413 10453
rect 24429 10389 24493 10453
rect 24509 10389 24573 10453
rect 24589 10389 24653 10453
rect 24669 10389 24733 10453
rect 24749 10389 24813 10453
rect 24829 10389 24893 10453
rect 24909 10389 24973 10453
rect 24989 10389 25053 10453
rect 25069 10389 25133 10453
rect 25149 10389 25213 10453
rect 25229 10389 25293 10453
rect 25309 10389 25373 10453
rect 25389 10389 25453 10453
rect 26309 10389 26373 10453
rect 26389 10389 26453 10453
rect 26469 10389 26533 10453
rect 26549 10389 26613 10453
rect 26629 10389 26693 10453
rect 26709 10389 26773 10453
rect 26789 10389 26853 10453
rect 26869 10389 26933 10453
rect 26949 10389 27013 10453
rect 27029 10389 27093 10453
rect 27109 10389 27173 10453
rect 27189 10389 27253 10453
rect 27269 10389 27333 10453
rect 27349 10389 27413 10453
rect 27429 10389 27493 10453
rect 27509 10389 27573 10453
rect 27589 10389 27653 10453
rect 27669 10389 27733 10453
rect 27749 10389 27813 10453
rect 27829 10389 27893 10453
rect 27909 10389 27973 10453
rect 27989 10389 28053 10453
rect 28069 10389 28133 10453
rect 28149 10389 28213 10453
rect 28229 10389 28293 10453
rect 28309 10389 28373 10453
rect 28389 10389 28453 10453
rect 28469 10389 28533 10453
rect 28549 10389 28613 10453
rect 28629 10389 28693 10453
rect 28709 10389 28773 10453
rect 28789 10389 28853 10453
rect 28869 10389 28933 10453
rect 28949 10389 29013 10453
rect 29029 10389 29093 10453
rect 29109 10389 29173 10453
rect 29189 10389 29253 10453
rect 29269 10389 29333 10453
rect 29349 10389 29413 10453
rect 29429 10389 29493 10453
rect 29509 10389 29573 10453
rect 29589 10389 29653 10453
rect 29669 10389 29733 10453
rect 29749 10389 29813 10453
rect 29829 10389 29893 10453
rect 29909 10389 29973 10453
rect 29989 10389 30053 10453
rect 30069 10389 30133 10453
rect 30149 10389 30213 10453
rect 30229 10389 30293 10453
rect 30309 10389 30373 10453
rect 30389 10389 30453 10453
rect 30469 10389 30533 10453
rect 30549 10389 30613 10453
rect 30629 10389 30693 10453
rect 30709 10389 30773 10453
rect 30789 10389 30853 10453
rect 30869 10389 30933 10453
rect 30949 10389 31013 10453
rect 31029 10389 31093 10453
rect 31109 10389 31173 10453
rect 31189 10389 31253 10453
rect 31269 10389 31333 10453
rect 31349 10389 31413 10453
rect 31429 10389 31493 10453
rect 31509 10389 31573 10453
rect 31589 10389 31653 10453
rect 31669 10389 31733 10453
rect 31749 10389 31813 10453
rect 31829 10389 31893 10453
rect 31909 10389 31973 10453
rect 31989 10389 32053 10453
rect 32069 10389 32133 10453
rect 32149 10389 32213 10453
rect 32229 10389 32293 10453
rect 32309 10389 32373 10453
rect 32389 10389 32453 10453
rect 21476 8895 21540 8910
rect 21476 8846 21478 8895
rect 21478 8846 21534 8895
rect 21534 8846 21540 8895
rect 21476 8759 21478 8800
rect 21478 8759 21534 8800
rect 21534 8759 21540 8800
rect 21476 8736 21540 8759
<< mimcap >>
rect -8619 16520 -2619 16568
rect -8619 10616 -8571 16520
rect -8274 16177 -8038 16413
rect -7954 16177 -7718 16413
rect -2667 10616 -2619 16520
rect -8619 10568 -2619 10616
rect -1619 16520 4381 16568
rect -1619 10616 -1571 16520
rect -1274 16177 -1038 16413
rect -954 16177 -718 16413
rect 4333 10616 4381 16520
rect -1619 10568 4381 10616
rect 5381 16520 11381 16568
rect 5381 10616 5429 16520
rect 5726 16177 5962 16413
rect 6046 16177 6282 16413
rect 11333 10616 11381 16520
rect 5381 10568 11381 10616
rect 12381 16520 18381 16568
rect 12381 10616 12429 16520
rect 12726 16177 12962 16413
rect 13046 16177 13282 16413
rect 18333 10616 18381 16520
rect 12381 10568 18381 10616
rect 19381 16520 25381 16568
rect 19381 10616 19429 16520
rect 19726 16177 19962 16413
rect 20046 16177 20282 16413
rect 25333 10616 25381 16520
rect 19381 10568 25381 10616
rect 26381 16520 32381 16568
rect 26381 10616 26429 16520
rect 26726 16177 26962 16413
rect 27046 16177 27282 16413
rect 32333 10616 32381 16520
rect 26381 10568 32381 10616
<< mimcapcontact >>
rect -8571 16413 -2667 16520
rect -8571 16177 -8274 16413
rect -8038 16177 -7954 16413
rect -7718 16177 -2667 16413
rect -8571 10616 -2667 16177
rect -1571 16413 4333 16520
rect -1571 16177 -1274 16413
rect -1038 16177 -954 16413
rect -718 16177 4333 16413
rect -1571 10616 4333 16177
rect 5429 16413 11333 16520
rect 5429 16177 5726 16413
rect 5962 16177 6046 16413
rect 6282 16177 11333 16413
rect 5429 10616 11333 16177
rect 12429 16413 18333 16520
rect 12429 16177 12726 16413
rect 12962 16177 13046 16413
rect 13282 16177 18333 16413
rect 12429 10616 18333 16177
rect 19429 16413 25333 16520
rect 19429 16177 19726 16413
rect 19962 16177 20046 16413
rect 20282 16177 25333 16413
rect 19429 10616 25333 16177
rect 26429 16413 32333 16520
rect 26429 16177 26726 16413
rect 26962 16177 27046 16413
rect 27282 16177 32333 16413
rect 26429 10616 32333 16177
<< metal4 >>
rect -8580 17163 32342 17218
rect -8580 16927 -8274 17163
rect -8038 16927 -7954 17163
rect -7718 16927 -1274 17163
rect -1038 16927 -954 17163
rect -718 16927 5726 17163
rect 5962 16927 6046 17163
rect 6282 17106 12726 17163
rect 6282 17042 11724 17106
rect 11788 17042 12726 17106
rect 6282 16996 12726 17042
rect 6282 16932 11724 16996
rect 11788 16932 12726 16996
rect 6282 16927 12726 16932
rect 12962 16927 13046 17163
rect 13282 16927 19726 17163
rect 19962 16927 20046 17163
rect 20282 16927 26726 17163
rect 26962 16927 27046 17163
rect 27282 16927 32342 17163
rect -8580 16873 32342 16927
rect -8580 16520 -2658 16529
rect -8580 10616 -8571 16520
rect -2667 10616 -2658 16520
rect -8580 10607 -2658 10616
rect -1580 16520 4342 16529
rect -1580 10616 -1571 16520
rect 4333 10616 4342 16520
rect -1580 10607 4342 10616
rect 5420 16520 11342 16529
rect 5420 10616 5429 16520
rect 11333 10616 11342 16520
rect 5420 10607 11342 10616
rect 12420 16520 18342 16529
rect 12420 10616 12429 16520
rect 18333 10616 18342 16520
rect 12420 10607 18342 10616
rect 19420 16520 25342 16529
rect 19420 10616 19429 16520
rect 25333 10616 25342 16520
rect 19420 10607 25342 10616
rect 26420 16520 32342 16529
rect 26420 10616 26429 16520
rect 32333 10616 32342 16520
rect 26420 10607 32342 10616
rect -8707 10453 -2531 10469
rect -8707 10389 -8691 10453
rect -8627 10389 -8611 10453
rect -8547 10389 -8531 10453
rect -8467 10389 -8451 10453
rect -8387 10389 -8371 10453
rect -8307 10389 -8291 10453
rect -8227 10389 -8211 10453
rect -8147 10389 -8131 10453
rect -8067 10389 -8051 10453
rect -7987 10389 -7971 10453
rect -7907 10389 -7891 10453
rect -7827 10389 -7811 10453
rect -7747 10389 -7731 10453
rect -7667 10389 -7651 10453
rect -7587 10389 -7571 10453
rect -7507 10389 -7491 10453
rect -7427 10389 -7411 10453
rect -7347 10389 -7331 10453
rect -7267 10389 -7251 10453
rect -7187 10389 -7171 10453
rect -7107 10389 -7091 10453
rect -7027 10389 -7011 10453
rect -6947 10389 -6931 10453
rect -6867 10389 -6851 10453
rect -6787 10389 -6771 10453
rect -6707 10389 -6691 10453
rect -6627 10389 -6611 10453
rect -6547 10389 -6531 10453
rect -6467 10389 -6451 10453
rect -6387 10389 -6371 10453
rect -6307 10389 -6291 10453
rect -6227 10389 -6211 10453
rect -6147 10389 -6131 10453
rect -6067 10389 -6051 10453
rect -5987 10389 -5971 10453
rect -5907 10389 -5891 10453
rect -5827 10389 -5811 10453
rect -5747 10389 -5731 10453
rect -5667 10389 -5651 10453
rect -5587 10389 -5571 10453
rect -5507 10389 -5491 10453
rect -5427 10389 -5411 10453
rect -5347 10389 -5331 10453
rect -5267 10389 -5251 10453
rect -5187 10389 -5171 10453
rect -5107 10389 -5091 10453
rect -5027 10389 -5011 10453
rect -4947 10389 -4931 10453
rect -4867 10389 -4851 10453
rect -4787 10389 -4771 10453
rect -4707 10389 -4691 10453
rect -4627 10389 -4611 10453
rect -4547 10389 -4531 10453
rect -4467 10389 -4451 10453
rect -4387 10389 -4371 10453
rect -4307 10389 -4291 10453
rect -4227 10389 -4211 10453
rect -4147 10389 -4131 10453
rect -4067 10389 -4051 10453
rect -3987 10389 -3971 10453
rect -3907 10389 -3891 10453
rect -3827 10389 -3811 10453
rect -3747 10389 -3731 10453
rect -3667 10389 -3651 10453
rect -3587 10389 -3571 10453
rect -3507 10389 -3491 10453
rect -3427 10389 -3411 10453
rect -3347 10389 -3331 10453
rect -3267 10389 -3251 10453
rect -3187 10389 -3171 10453
rect -3107 10389 -3091 10453
rect -3027 10389 -3011 10453
rect -2947 10389 -2931 10453
rect -2867 10389 -2851 10453
rect -2787 10389 -2771 10453
rect -2707 10389 -2691 10453
rect -2627 10389 -2611 10453
rect -2547 10389 -2531 10453
rect -8707 10373 -2531 10389
rect -1707 10453 4469 10469
rect -1707 10389 -1691 10453
rect -1627 10389 -1611 10453
rect -1547 10389 -1531 10453
rect -1467 10389 -1451 10453
rect -1387 10389 -1371 10453
rect -1307 10389 -1291 10453
rect -1227 10389 -1211 10453
rect -1147 10389 -1131 10453
rect -1067 10389 -1051 10453
rect -987 10389 -971 10453
rect -907 10389 -891 10453
rect -827 10389 -811 10453
rect -747 10389 -731 10453
rect -667 10389 -651 10453
rect -587 10389 -571 10453
rect -507 10389 -491 10453
rect -427 10389 -411 10453
rect -347 10389 -331 10453
rect -267 10389 -251 10453
rect -187 10389 -171 10453
rect -107 10389 -91 10453
rect -27 10389 -11 10453
rect 53 10389 69 10453
rect 133 10389 149 10453
rect 213 10389 229 10453
rect 293 10389 309 10453
rect 373 10389 389 10453
rect 453 10389 469 10453
rect 533 10389 549 10453
rect 613 10389 629 10453
rect 693 10389 709 10453
rect 773 10389 789 10453
rect 853 10389 869 10453
rect 933 10389 949 10453
rect 1013 10389 1029 10453
rect 1093 10389 1109 10453
rect 1173 10389 1189 10453
rect 1253 10389 1269 10453
rect 1333 10389 1349 10453
rect 1413 10389 1429 10453
rect 1493 10389 1509 10453
rect 1573 10389 1589 10453
rect 1653 10389 1669 10453
rect 1733 10389 1749 10453
rect 1813 10389 1829 10453
rect 1893 10389 1909 10453
rect 1973 10389 1989 10453
rect 2053 10389 2069 10453
rect 2133 10389 2149 10453
rect 2213 10389 2229 10453
rect 2293 10389 2309 10453
rect 2373 10389 2389 10453
rect 2453 10389 2469 10453
rect 2533 10389 2549 10453
rect 2613 10389 2629 10453
rect 2693 10389 2709 10453
rect 2773 10389 2789 10453
rect 2853 10389 2869 10453
rect 2933 10389 2949 10453
rect 3013 10389 3029 10453
rect 3093 10389 3109 10453
rect 3173 10389 3189 10453
rect 3253 10389 3269 10453
rect 3333 10389 3349 10453
rect 3413 10389 3429 10453
rect 3493 10389 3509 10453
rect 3573 10389 3589 10453
rect 3653 10389 3669 10453
rect 3733 10389 3749 10453
rect 3813 10389 3829 10453
rect 3893 10389 3909 10453
rect 3973 10389 3989 10453
rect 4053 10389 4069 10453
rect 4133 10389 4149 10453
rect 4213 10389 4229 10453
rect 4293 10389 4309 10453
rect 4373 10389 4389 10453
rect 4453 10389 4469 10453
rect -1707 10373 4469 10389
rect 5293 10453 11469 10469
rect 5293 10389 5309 10453
rect 5373 10389 5389 10453
rect 5453 10389 5469 10453
rect 5533 10389 5549 10453
rect 5613 10389 5629 10453
rect 5693 10389 5709 10453
rect 5773 10389 5789 10453
rect 5853 10389 5869 10453
rect 5933 10389 5949 10453
rect 6013 10389 6029 10453
rect 6093 10389 6109 10453
rect 6173 10389 6189 10453
rect 6253 10389 6269 10453
rect 6333 10389 6349 10453
rect 6413 10389 6429 10453
rect 6493 10389 6509 10453
rect 6573 10389 6589 10453
rect 6653 10389 6669 10453
rect 6733 10389 6749 10453
rect 6813 10389 6829 10453
rect 6893 10389 6909 10453
rect 6973 10389 6989 10453
rect 7053 10389 7069 10453
rect 7133 10389 7149 10453
rect 7213 10389 7229 10453
rect 7293 10389 7309 10453
rect 7373 10389 7389 10453
rect 7453 10389 7469 10453
rect 7533 10389 7549 10453
rect 7613 10389 7629 10453
rect 7693 10389 7709 10453
rect 7773 10389 7789 10453
rect 7853 10389 7869 10453
rect 7933 10389 7949 10453
rect 8013 10389 8029 10453
rect 8093 10389 8109 10453
rect 8173 10389 8189 10453
rect 8253 10389 8269 10453
rect 8333 10389 8349 10453
rect 8413 10389 8429 10453
rect 8493 10389 8509 10453
rect 8573 10389 8589 10453
rect 8653 10389 8669 10453
rect 8733 10389 8749 10453
rect 8813 10389 8829 10453
rect 8893 10389 8909 10453
rect 8973 10389 8989 10453
rect 9053 10389 9069 10453
rect 9133 10389 9149 10453
rect 9213 10389 9229 10453
rect 9293 10389 9309 10453
rect 9373 10389 9389 10453
rect 9453 10389 9469 10453
rect 9533 10389 9549 10453
rect 9613 10389 9629 10453
rect 9693 10389 9709 10453
rect 9773 10389 9789 10453
rect 9853 10389 9869 10453
rect 9933 10389 9949 10453
rect 10013 10389 10029 10453
rect 10093 10389 10109 10453
rect 10173 10389 10189 10453
rect 10253 10389 10269 10453
rect 10333 10389 10349 10453
rect 10413 10389 10429 10453
rect 10493 10389 10509 10453
rect 10573 10389 10589 10453
rect 10653 10389 10669 10453
rect 10733 10389 10749 10453
rect 10813 10389 10829 10453
rect 10893 10389 10909 10453
rect 10973 10389 10989 10453
rect 11053 10389 11069 10453
rect 11133 10389 11149 10453
rect 11213 10389 11229 10453
rect 11293 10389 11309 10453
rect 11373 10389 11389 10453
rect 11453 10389 11469 10453
rect 5293 10373 11469 10389
rect 12293 10453 18469 10469
rect 12293 10389 12309 10453
rect 12373 10389 12389 10453
rect 12453 10389 12469 10453
rect 12533 10389 12549 10453
rect 12613 10389 12629 10453
rect 12693 10389 12709 10453
rect 12773 10389 12789 10453
rect 12853 10389 12869 10453
rect 12933 10389 12949 10453
rect 13013 10389 13029 10453
rect 13093 10389 13109 10453
rect 13173 10389 13189 10453
rect 13253 10389 13269 10453
rect 13333 10389 13349 10453
rect 13413 10389 13429 10453
rect 13493 10389 13509 10453
rect 13573 10389 13589 10453
rect 13653 10389 13669 10453
rect 13733 10389 13749 10453
rect 13813 10389 13829 10453
rect 13893 10389 13909 10453
rect 13973 10389 13989 10453
rect 14053 10389 14069 10453
rect 14133 10389 14149 10453
rect 14213 10389 14229 10453
rect 14293 10389 14309 10453
rect 14373 10389 14389 10453
rect 14453 10389 14469 10453
rect 14533 10389 14549 10453
rect 14613 10389 14629 10453
rect 14693 10389 14709 10453
rect 14773 10389 14789 10453
rect 14853 10389 14869 10453
rect 14933 10389 14949 10453
rect 15013 10389 15029 10453
rect 15093 10389 15109 10453
rect 15173 10389 15189 10453
rect 15253 10389 15269 10453
rect 15333 10389 15349 10453
rect 15413 10389 15429 10453
rect 15493 10389 15509 10453
rect 15573 10389 15589 10453
rect 15653 10389 15669 10453
rect 15733 10389 15749 10453
rect 15813 10389 15829 10453
rect 15893 10389 15909 10453
rect 15973 10389 15989 10453
rect 16053 10389 16069 10453
rect 16133 10389 16149 10453
rect 16213 10389 16229 10453
rect 16293 10389 16309 10453
rect 16373 10389 16389 10453
rect 16453 10389 16469 10453
rect 16533 10389 16549 10453
rect 16613 10389 16629 10453
rect 16693 10389 16709 10453
rect 16773 10389 16789 10453
rect 16853 10389 16869 10453
rect 16933 10389 16949 10453
rect 17013 10389 17029 10453
rect 17093 10389 17109 10453
rect 17173 10389 17189 10453
rect 17253 10389 17269 10453
rect 17333 10389 17349 10453
rect 17413 10389 17429 10453
rect 17493 10389 17509 10453
rect 17573 10389 17589 10453
rect 17653 10389 17669 10453
rect 17733 10389 17749 10453
rect 17813 10389 17829 10453
rect 17893 10389 17909 10453
rect 17973 10389 17989 10453
rect 18053 10389 18069 10453
rect 18133 10389 18149 10453
rect 18213 10389 18229 10453
rect 18293 10389 18309 10453
rect 18373 10389 18389 10453
rect 18453 10389 18469 10453
rect 12293 10373 18469 10389
rect 19293 10453 25469 10469
rect 19293 10389 19309 10453
rect 19373 10389 19389 10453
rect 19453 10389 19469 10453
rect 19533 10389 19549 10453
rect 19613 10389 19629 10453
rect 19693 10389 19709 10453
rect 19773 10389 19789 10453
rect 19853 10389 19869 10453
rect 19933 10389 19949 10453
rect 20013 10389 20029 10453
rect 20093 10389 20109 10453
rect 20173 10389 20189 10453
rect 20253 10389 20269 10453
rect 20333 10389 20349 10453
rect 20413 10389 20429 10453
rect 20493 10389 20509 10453
rect 20573 10389 20589 10453
rect 20653 10389 20669 10453
rect 20733 10389 20749 10453
rect 20813 10389 20829 10453
rect 20893 10389 20909 10453
rect 20973 10389 20989 10453
rect 21053 10389 21069 10453
rect 21133 10389 21149 10453
rect 21213 10389 21229 10453
rect 21293 10389 21309 10453
rect 21373 10389 21389 10453
rect 21453 10389 21469 10453
rect 21533 10389 21549 10453
rect 21613 10389 21629 10453
rect 21693 10389 21709 10453
rect 21773 10389 21789 10453
rect 21853 10389 21869 10453
rect 21933 10389 21949 10453
rect 22013 10389 22029 10453
rect 22093 10389 22109 10453
rect 22173 10389 22189 10453
rect 22253 10389 22269 10453
rect 22333 10389 22349 10453
rect 22413 10389 22429 10453
rect 22493 10389 22509 10453
rect 22573 10389 22589 10453
rect 22653 10389 22669 10453
rect 22733 10389 22749 10453
rect 22813 10389 22829 10453
rect 22893 10389 22909 10453
rect 22973 10389 22989 10453
rect 23053 10389 23069 10453
rect 23133 10389 23149 10453
rect 23213 10389 23229 10453
rect 23293 10389 23309 10453
rect 23373 10389 23389 10453
rect 23453 10389 23469 10453
rect 23533 10389 23549 10453
rect 23613 10389 23629 10453
rect 23693 10389 23709 10453
rect 23773 10389 23789 10453
rect 23853 10389 23869 10453
rect 23933 10389 23949 10453
rect 24013 10389 24029 10453
rect 24093 10389 24109 10453
rect 24173 10389 24189 10453
rect 24253 10389 24269 10453
rect 24333 10389 24349 10453
rect 24413 10389 24429 10453
rect 24493 10389 24509 10453
rect 24573 10389 24589 10453
rect 24653 10389 24669 10453
rect 24733 10389 24749 10453
rect 24813 10389 24829 10453
rect 24893 10389 24909 10453
rect 24973 10389 24989 10453
rect 25053 10389 25069 10453
rect 25133 10389 25149 10453
rect 25213 10389 25229 10453
rect 25293 10389 25309 10453
rect 25373 10389 25389 10453
rect 25453 10389 25469 10453
rect 19293 10373 25469 10389
rect 26293 10453 32469 10469
rect 26293 10389 26309 10453
rect 26373 10389 26389 10453
rect 26453 10389 26469 10453
rect 26533 10389 26549 10453
rect 26613 10389 26629 10453
rect 26693 10389 26709 10453
rect 26773 10389 26789 10453
rect 26853 10389 26869 10453
rect 26933 10389 26949 10453
rect 27013 10389 27029 10453
rect 27093 10389 27109 10453
rect 27173 10389 27189 10453
rect 27253 10389 27269 10453
rect 27333 10389 27349 10453
rect 27413 10389 27429 10453
rect 27493 10389 27509 10453
rect 27573 10389 27589 10453
rect 27653 10389 27669 10453
rect 27733 10389 27749 10453
rect 27813 10389 27829 10453
rect 27893 10389 27909 10453
rect 27973 10389 27989 10453
rect 28053 10389 28069 10453
rect 28133 10389 28149 10453
rect 28213 10389 28229 10453
rect 28293 10389 28309 10453
rect 28373 10389 28389 10453
rect 28453 10389 28469 10453
rect 28533 10389 28549 10453
rect 28613 10389 28629 10453
rect 28693 10389 28709 10453
rect 28773 10389 28789 10453
rect 28853 10389 28869 10453
rect 28933 10389 28949 10453
rect 29013 10389 29029 10453
rect 29093 10389 29109 10453
rect 29173 10389 29189 10453
rect 29253 10389 29269 10453
rect 29333 10389 29349 10453
rect 29413 10389 29429 10453
rect 29493 10389 29509 10453
rect 29573 10389 29589 10453
rect 29653 10389 29669 10453
rect 29733 10389 29749 10453
rect 29813 10389 29829 10453
rect 29893 10389 29909 10453
rect 29973 10389 29989 10453
rect 30053 10389 30069 10453
rect 30133 10389 30149 10453
rect 30213 10389 30229 10453
rect 30293 10389 30309 10453
rect 30373 10389 30389 10453
rect 30453 10389 30469 10453
rect 30533 10389 30549 10453
rect 30613 10389 30629 10453
rect 30693 10389 30709 10453
rect 30773 10389 30789 10453
rect 30853 10389 30869 10453
rect 30933 10389 30949 10453
rect 31013 10389 31029 10453
rect 31093 10389 31109 10453
rect 31173 10389 31189 10453
rect 31253 10389 31269 10453
rect 31333 10389 31349 10453
rect 31413 10389 31429 10453
rect 31493 10389 31509 10453
rect 31573 10389 31589 10453
rect 31653 10389 31669 10453
rect 31733 10389 31749 10453
rect 31813 10389 31829 10453
rect 31893 10389 31909 10453
rect 31973 10389 31989 10453
rect 32053 10389 32069 10453
rect 32133 10389 32149 10453
rect 32213 10389 32229 10453
rect 32293 10389 32309 10453
rect 32373 10389 32389 10453
rect 32453 10389 32469 10453
rect 26293 10373 32469 10389
rect -8707 10181 32469 10373
rect 21470 8910 21546 10181
rect 21470 8846 21476 8910
rect 21540 8846 21546 8910
rect 21470 8800 21546 8846
rect 21470 8736 21476 8800
rect 21540 8736 21546 8800
rect 21470 8730 21546 8736
<< via4 >>
rect -8274 16927 -8038 17163
rect -7954 16927 -7718 17163
rect -1274 16927 -1038 17163
rect -954 16927 -718 17163
rect 5726 16927 5962 17163
rect 6046 16927 6282 17163
rect 12726 16927 12962 17163
rect 13046 16927 13282 17163
rect 19726 16927 19962 17163
rect 20046 16927 20282 17163
rect 26726 16927 26962 17163
rect 27046 16927 27282 17163
rect -8274 16177 -8038 16413
rect -7954 16177 -7718 16413
rect -1274 16177 -1038 16413
rect -954 16177 -718 16413
rect 5726 16177 5962 16413
rect 6046 16177 6282 16413
rect 12726 16177 12962 16413
rect 13046 16177 13282 16413
rect 19726 16177 19962 16413
rect 20046 16177 20282 16413
rect 26726 16177 26962 16413
rect 27046 16177 27282 16413
<< metal5 >>
rect -8298 17163 -7694 17187
rect -8298 16927 -8274 17163
rect -8038 16927 -7954 17163
rect -7718 16927 -7694 17163
rect -8298 16413 -7694 16927
rect -8298 16177 -8274 16413
rect -8038 16177 -7954 16413
rect -7718 16177 -7694 16413
rect -8298 16153 -7694 16177
rect -1298 17163 -694 17187
rect -1298 16927 -1274 17163
rect -1038 16927 -954 17163
rect -718 16927 -694 17163
rect -1298 16413 -694 16927
rect -1298 16177 -1274 16413
rect -1038 16177 -954 16413
rect -718 16177 -694 16413
rect -1298 16153 -694 16177
rect 5702 17163 6306 17187
rect 5702 16927 5726 17163
rect 5962 16927 6046 17163
rect 6282 16927 6306 17163
rect 5702 16413 6306 16927
rect 5702 16177 5726 16413
rect 5962 16177 6046 16413
rect 6282 16177 6306 16413
rect 5702 16153 6306 16177
rect 12702 17163 13306 17187
rect 12702 16927 12726 17163
rect 12962 16927 13046 17163
rect 13282 16927 13306 17163
rect 12702 16413 13306 16927
rect 12702 16177 12726 16413
rect 12962 16177 13046 16413
rect 13282 16177 13306 16413
rect 12702 16153 13306 16177
rect 19702 17163 20306 17187
rect 19702 16927 19726 17163
rect 19962 16927 20046 17163
rect 20282 16927 20306 17163
rect 19702 16413 20306 16927
rect 19702 16177 19726 16413
rect 19962 16177 20046 16413
rect 20282 16177 20306 16413
rect 19702 16153 20306 16177
rect 26702 17163 27306 17187
rect 26702 16927 26726 17163
rect 26962 16927 27046 17163
rect 27282 16927 27306 17163
rect 26702 16413 27306 16927
rect 26702 16177 26726 16413
rect 26962 16177 27046 16413
rect 27282 16177 27306 16413
rect 26702 16153 27306 16177
<< labels >>
flabel metal2 s -9198 3414 -9048 3498 2 FreeSans 2000 0 0 0 in_n
port 5 nsew
flabel metal2 s 33680 3414 33850 3498 2 FreeSans 2000 0 0 0 in_p
port 6 nsew
rlabel metal1 -9200 8950 -9080 9070 1 vdd
port 7 n
rlabel metal1 -9200 2280 -9070 2420 1 bias
port 8 n
rlabel metal1 33530 3730 33850 3980 1 out
port 9 n
rlabel metal1 -9200 490 -8990 720 1 vss
port 10 n
<< properties >>
string FIXED_BBOX 26281 10468 32481 16668
<< end >>
