magic
tech sky130A
timestamp 1635946216
<< error_p >>
rect 69 1063 70 1080
rect 87 1063 89 1080
rect 6 1011 23 1012
rect 135 1011 152 1012
rect 6 1003 23 1004
rect 135 1003 152 1004
rect 6 984 23 985
rect 135 984 152 985
rect 6 977 23 978
rect 135 977 152 978
rect 6 967 23 968
rect 135 967 152 968
rect 6 948 23 949
rect 135 948 152 949
rect 6 943 23 944
rect 135 943 152 944
rect 6 931 23 932
rect 135 931 152 932
rect 6 912 23 913
rect 135 912 152 913
rect 6 909 23 910
rect 135 909 152 910
rect 6 895 23 896
rect 135 895 152 896
rect 6 875 23 877
rect 135 875 152 877
rect 6 859 23 860
rect 135 859 152 860
rect 6 840 23 842
rect 135 840 152 842
rect 6 823 23 824
rect 135 823 152 824
rect 6 807 23 808
rect 135 807 152 808
rect 6 804 23 805
rect 135 804 152 805
rect 6 787 23 788
rect 135 787 152 788
rect 6 773 23 774
rect 135 773 152 774
rect 6 768 23 769
rect 135 768 152 769
rect 6 751 23 752
rect 135 751 152 752
rect 6 739 23 740
rect 135 739 152 740
rect 6 732 23 733
rect 135 732 152 733
rect 6 715 23 716
rect 135 715 152 716
rect 6 705 23 706
rect 135 705 152 706
rect 6 696 23 697
rect 135 696 152 697
rect 6 679 23 680
rect 135 679 152 680
rect 6 671 23 672
rect 135 671 152 672
rect 6 660 23 661
rect 135 660 152 661
rect 6 643 23 644
rect 135 643 152 644
rect 6 637 23 638
rect 135 637 152 638
rect 6 624 23 625
rect 135 624 152 625
rect 6 607 23 608
rect 135 607 152 608
rect 6 603 23 604
rect 135 603 152 604
rect 6 588 23 589
rect 135 588 152 589
rect 6 571 23 572
rect 135 571 152 572
rect 6 569 23 570
rect 135 569 152 570
rect 6 552 23 553
rect 135 552 152 553
rect 6 535 23 536
rect 135 535 152 536
rect 6 516 23 517
rect 135 516 152 517
rect 6 501 23 502
rect 135 501 152 502
rect 6 499 23 500
rect 135 499 152 500
rect 6 480 23 481
rect 135 480 152 481
rect 6 467 23 468
rect 135 467 152 468
rect 6 463 23 464
rect 135 463 152 464
rect 6 444 23 445
rect 135 444 152 445
rect 6 433 23 434
rect 135 433 152 434
rect 6 427 23 428
rect 135 427 152 428
rect 6 408 23 409
rect 135 408 152 409
rect 6 399 23 400
rect 135 399 152 400
rect 6 391 23 392
rect 135 391 152 392
rect 6 372 23 373
rect 135 372 152 373
rect 6 365 23 366
rect 135 365 152 366
rect 6 355 23 356
rect 135 355 152 356
rect 6 336 23 337
rect 135 336 152 337
rect 6 331 23 332
rect 135 331 152 332
rect 6 319 23 320
rect 135 319 152 320
rect 6 300 23 301
rect 135 300 152 301
rect 6 297 23 298
rect 135 297 152 298
rect 6 283 23 284
rect 135 283 152 284
rect 6 263 23 265
rect 135 263 152 265
rect 6 247 23 248
rect 135 247 152 248
rect 6 228 23 230
rect 135 228 152 230
rect 6 211 23 212
rect 135 211 152 212
rect 6 195 23 196
rect 135 195 152 196
rect 6 192 23 193
rect 135 192 152 193
rect 6 175 23 176
rect 135 175 152 176
rect 6 161 23 162
rect 135 161 152 162
rect 6 156 23 157
rect 135 156 152 157
rect 6 139 23 140
rect 135 139 152 140
rect 6 127 23 128
rect 135 127 152 128
rect 6 120 23 121
rect 135 120 152 121
rect 6 103 23 104
rect 135 103 152 104
rect 6 93 23 94
rect 135 93 152 94
rect 6 84 23 85
rect 135 84 152 85
rect 69 8 70 25
rect 87 8 89 25
use sky130_fd_pr__nfet_g5v0d10v5_9A4VCP  sky130_fd_pr__nfet_g5v0d10v5_9A4VCP_0
timestamp 1635946216
transform 1 0 79 0 1 544
box -92 -544 92 544
<< end >>
