* SPICE3 file created from /mnt/c/Users/Harry/magic-practice/caravel_user_project_analog/comparator/decision.ext - technology: sky130A

.option scale=1u

X0 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=-0 pd=0 as=-0 ps=0 w=1.5e+06 l=500000
X1 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=-0 pd=0 as=-0 ps=0 w=1.5e+06 l=500000
X2 VOP VPAMP VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=-0 ps=0 w=1.5e+06 l=500000
X3 VON VNAMP VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=-0 ps=0 w=1.5e+06 l=500000
X4 ISINK VOP VOP VGND sky130_fd_pr__nfet_03v3_nvt ad=-0 pd=0 as=0 ps=0 w=1e+06 l=600000
X5 VGND VGND VGND VGND sky130_fd_pr__nfet_03v3_nvt ad=-0 pd=0 as=-0 ps=0 w=1e+06 l=600000
X6 ISINK VON VON VGND sky130_fd_pr__nfet_03v3_nvt ad=-0 pd=0 as=0 ps=0 w=1e+06 l=600000
X7 ISINK VOP VON VGND sky130_fd_pr__nfet_03v3_nvt ad=-0 pd=0 as=0 ps=0 w=1e+06 l=600000
X8 ISINK VON VOP VGND sky130_fd_pr__nfet_03v3_nvt ad=-0 pd=0 as=0 ps=0 w=1e+06 l=600000
X9 VGND VGND VGND VGND sky130_fd_pr__nfet_03v3_nvt ad=-0 pd=0 as=-0 ps=0 w=1e+06 l=600000
X10 VGND ISINK ISINK VGND sky130_fd_pr__nfet_03v3_nvt ad=-0 pd=0 as=-0 ps=0 w=1e+06 l=600000
X11 VGND VGND VGND VGND sky130_fd_pr__nfet_03v3_nvt ad=-0 pd=0 as=-0 ps=0 w=1e+06 l=600000
X12 VGND VGND VGND VGND sky130_fd_pr__nfet_03v3_nvt ad=-0 pd=0 as=-0 ps=0 w=1e+06 l=600000
C0 VPWR VGND 6.67fF
C1 ISINK VGND 2.29fF
C2 VON VGND 2.41fF
