* NGSPICE file created from preamp.ext - technology: sky130A

X0 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=-0p pd=0u as=-0p ps=0u w=1.5e+06u l=500000u
X1 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=-0p pd=0u as=-0p ps=0u w=1.5e+06u l=500000u
X2 VPAMP VPAMP VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=-0p ps=0u w=1.5e+06u l=500000u
X3 VNAMP VNAMP VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=-0p ps=0u w=1.5e+06u l=500000u
X4 VGND BIASN VI VGND sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=-0p ps=0u w=1e+06u l=600000u
X5 VGND VGND VGND VGND sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=600000u
X6 VI BIASN VGND VGND sky130_fd_pr__nfet_03v3_nvt ad=-0p pd=0u as=0p ps=0u w=1e+06u l=600000u
X7 VGND VGND VGND VGND sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=600000u
X8 VGND VGND VGND VGND sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=600000u
X9 VGND VGND VGND VGND sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=600000u
X10 VGND VGND VGND VGND sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=600000u
X11 VGND VGND VGND VGND sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=600000u
X12 VI VN VNAMP VGND sky130_fd_pr__nfet_03v3_nvt ad=-0p pd=0u as=-0p ps=0u w=1e+06u l=600000u
X13 VI VP VPAMP VGND sky130_fd_pr__nfet_03v3_nvt ad=-0p pd=0u as=-0p ps=0u w=1e+06u l=600000u
C0 VPWR VGND 8.16fF
