magic
tech sky130A
timestamp 1632928825
<< nwell >>
rect 210 -330 730 240
rect 930 -770 1320 -140
<< pwell >>
rect -250 -190 140 230
rect -310 -240 140 -190
rect -250 -270 140 -240
rect -250 -1040 -230 -270
rect -215 -1025 -115 -285
rect -110 -440 140 -270
rect -110 -1040 510 -440
rect -250 -1060 510 -1040
<< nmos >>
rect 280 -810 298 -710
rect 350 -810 368 -710
rect 60 -960 78 -860
rect 190 -1030 205 -930
<< pmos >>
rect 990 -460 1008 -160
rect 1060 -460 1078 -160
rect 990 -750 1005 -550
<< mvnmos >>
rect 20 110 120 170
rect 20 0 120 60
rect 20 -190 120 -130
rect 20 -300 120 -240
rect 60 -560 120 -460
rect 170 -560 230 -460
rect 280 -560 340 -460
rect 390 -560 450 -460
rect 60 -760 120 -660
<< mvpmos >>
rect 250 110 400 160
rect 250 10 400 60
rect 250 -150 400 -100
rect 250 -250 400 -200
<< ndiff >>
rect 240 -720 280 -710
rect 240 -800 250 -720
rect 270 -800 280 -720
rect 240 -810 280 -800
rect 298 -720 350 -710
rect 298 -800 310 -720
rect 340 -800 350 -720
rect 298 -810 350 -800
rect 368 -720 410 -710
rect 368 -800 380 -720
rect 400 -800 410 -720
rect 368 -810 410 -800
rect 20 -870 60 -860
rect 20 -950 30 -870
rect 50 -950 60 -870
rect 20 -960 60 -950
rect 78 -870 120 -860
rect 78 -950 90 -870
rect 110 -950 120 -870
rect 78 -960 120 -950
rect 150 -940 190 -930
rect 150 -1020 160 -940
rect 180 -1020 190 -940
rect 150 -1030 190 -1020
rect 205 -940 250 -930
rect 205 -1020 220 -940
rect 240 -1020 250 -940
rect 205 -1030 250 -1020
<< pdiff >>
rect 950 -170 990 -160
rect 950 -450 960 -170
rect 980 -450 990 -170
rect 950 -460 990 -450
rect 1008 -170 1060 -160
rect 1008 -450 1020 -170
rect 1050 -450 1060 -170
rect 1008 -460 1060 -450
rect 1078 -170 1120 -160
rect 1078 -450 1090 -170
rect 1110 -450 1120 -170
rect 1078 -460 1120 -450
rect 950 -560 990 -550
rect 950 -740 960 -560
rect 980 -740 990 -560
rect 950 -750 990 -740
rect 1005 -560 1050 -550
rect 1005 -740 1020 -560
rect 1040 -740 1050 -560
rect 1005 -750 1050 -740
<< mvndiff >>
rect 20 200 120 210
rect 20 180 30 200
rect 110 180 120 200
rect 20 170 120 180
rect 20 100 120 110
rect 20 70 30 100
rect 110 70 120 100
rect 20 60 120 70
rect 20 -10 120 0
rect 20 -30 30 -10
rect 110 -30 120 -10
rect 20 -40 120 -30
rect 20 -100 120 -90
rect 20 -120 30 -100
rect 110 -120 120 -100
rect 20 -130 120 -120
rect 20 -200 120 -190
rect 20 -230 30 -200
rect 110 -230 120 -200
rect 20 -240 120 -230
rect 20 -310 120 -300
rect 20 -330 30 -310
rect 110 -330 120 -310
rect 20 -340 120 -330
rect 20 -470 60 -460
rect 20 -550 30 -470
rect 50 -550 60 -470
rect 20 -560 60 -550
rect 120 -470 170 -460
rect 120 -550 130 -470
rect 160 -550 170 -470
rect 120 -560 170 -550
rect 230 -470 280 -460
rect 230 -550 240 -470
rect 270 -550 280 -470
rect 230 -560 280 -550
rect 340 -470 390 -460
rect 340 -550 350 -470
rect 380 -550 390 -470
rect 340 -560 390 -550
rect 450 -470 490 -460
rect 450 -550 460 -470
rect 480 -550 490 -470
rect 450 -560 490 -550
rect 20 -670 60 -660
rect 20 -750 30 -670
rect 50 -750 60 -670
rect 20 -760 60 -750
rect 120 -670 160 -660
rect 120 -750 130 -670
rect 150 -750 160 -670
rect 120 -760 160 -750
<< mvpdiff >>
rect 250 190 400 200
rect 250 170 260 190
rect 390 170 400 190
rect 250 160 400 170
rect 250 100 400 110
rect 250 70 260 100
rect 390 70 400 100
rect 250 60 400 70
rect 250 0 400 10
rect 250 -20 260 0
rect 390 -20 400 0
rect 250 -30 400 -20
rect 250 -70 400 -60
rect 250 -90 260 -70
rect 390 -90 400 -70
rect 250 -100 400 -90
rect 250 -160 400 -150
rect 250 -190 260 -160
rect 390 -190 400 -160
rect 250 -200 400 -190
rect 250 -260 400 -250
rect 250 -280 260 -260
rect 390 -280 400 -260
rect 250 -290 400 -280
<< ndiffc >>
rect 250 -800 270 -720
rect 310 -800 340 -720
rect 380 -800 400 -720
rect 30 -950 50 -870
rect 90 -950 110 -870
rect 160 -1020 180 -940
rect 220 -1020 240 -940
<< pdiffc >>
rect 960 -450 980 -170
rect 1020 -450 1050 -170
rect 1090 -450 1110 -170
rect 960 -740 980 -560
rect 1020 -740 1040 -560
<< mvndiffc >>
rect 30 180 110 200
rect 30 70 110 100
rect 30 -30 110 -10
rect 30 -120 110 -100
rect 30 -230 110 -200
rect 30 -330 110 -310
rect 30 -550 50 -470
rect 130 -550 160 -470
rect 240 -550 270 -470
rect 350 -550 380 -470
rect 460 -550 480 -470
rect 30 -750 50 -670
rect 130 -750 150 -670
<< mvpdiffc >>
rect 260 170 390 190
rect 260 70 390 100
rect 260 -20 390 0
rect 260 -90 390 -70
rect 260 -190 390 -160
rect 260 -280 390 -260
<< psubdiff >>
rect -230 -160 -215 -40
rect -115 -160 -100 -40
rect -230 -285 -100 -270
rect -230 -1025 -215 -285
rect -115 -1025 -100 -285
rect -230 -1040 -100 -1025
<< nsubdiff >>
rect 600 185 690 200
rect 600 -275 615 185
rect 600 -290 690 -275
rect 1200 -175 1300 -160
rect 1200 -735 1215 -175
rect 1285 -735 1300 -175
rect 1200 -750 1300 -735
<< psubdiffcont >>
rect -215 -160 -115 -40
rect -215 -1025 -115 -285
<< nsubdiffcont >>
rect 615 -275 690 185
rect 1215 -735 1285 -175
<< poly >>
rect -60 160 20 170
rect -60 120 -50 160
rect -10 120 20 160
rect -60 110 20 120
rect 120 110 150 170
rect 220 110 250 160
rect 400 150 550 160
rect 400 130 440 150
rect 460 130 550 150
rect 400 110 550 130
rect -60 50 20 60
rect -60 10 -50 50
rect -10 10 20 50
rect -60 0 20 10
rect 120 0 150 60
rect 220 10 250 60
rect 400 40 470 60
rect 400 20 440 40
rect 460 20 470 40
rect 400 10 470 20
rect 420 -100 470 10
rect -50 -190 20 -130
rect 120 -190 150 -130
rect 220 -150 250 -100
rect 400 -150 470 -100
rect -50 -200 0 -190
rect -50 -230 -40 -200
rect -10 -230 0 -200
rect -50 -240 0 -230
rect 500 -200 550 110
rect -50 -300 20 -240
rect 120 -300 150 -240
rect 220 -250 250 -200
rect 400 -250 550 -200
rect 990 -110 1030 -100
rect 990 -130 1000 -110
rect 1020 -130 1078 -110
rect 990 -140 1078 -130
rect 990 -160 1008 -140
rect 1060 -160 1078 -140
rect 160 -360 210 -350
rect 160 -370 170 -360
rect 60 -390 170 -370
rect 200 -370 210 -360
rect 200 -390 450 -370
rect 60 -400 450 -390
rect 60 -460 120 -400
rect 170 -460 230 -430
rect 280 -460 340 -430
rect 390 -460 450 -400
rect 990 -490 1008 -460
rect 1060 -490 1078 -460
rect 990 -550 1005 -520
rect 60 -590 120 -560
rect 170 -590 230 -560
rect 280 -580 340 -560
rect 280 -590 300 -580
rect -10 -610 30 -600
rect -10 -630 0 -610
rect 20 -620 30 -610
rect 170 -610 300 -590
rect 330 -610 340 -580
rect 390 -590 450 -560
rect 170 -620 340 -610
rect 20 -630 120 -620
rect -10 -640 120 -630
rect 60 -660 120 -640
rect 250 -660 310 -650
rect 250 -680 260 -660
rect 280 -680 310 -660
rect 250 -690 310 -680
rect 350 -660 395 -650
rect 350 -680 365 -660
rect 385 -680 395 -660
rect 350 -690 395 -680
rect 280 -710 298 -690
rect 350 -710 368 -690
rect 60 -790 120 -760
rect 440 -780 480 -770
rect 990 -780 1005 -750
rect 440 -800 450 -780
rect 470 -800 480 -780
rect 140 -820 180 -810
rect 60 -840 150 -820
rect 170 -840 180 -820
rect 280 -840 298 -810
rect 350 -840 368 -810
rect 60 -860 78 -840
rect 140 -850 180 -840
rect 440 -880 480 -800
rect 730 -790 1130 -780
rect 730 -830 740 -790
rect 840 -830 1020 -790
rect 1120 -830 1130 -790
rect 730 -840 1130 -830
rect 190 -910 480 -880
rect 190 -930 205 -910
rect 60 -990 78 -960
rect 190 -1060 205 -1030
<< polycont >>
rect -50 120 -10 160
rect 440 130 460 150
rect -50 10 -10 50
rect 440 20 460 40
rect -40 -230 -10 -200
rect 1000 -130 1020 -110
rect 170 -390 200 -360
rect 0 -630 20 -610
rect 300 -610 330 -580
rect 260 -680 280 -660
rect 365 -680 385 -660
rect 450 -800 470 -780
rect 150 -840 170 -820
rect 740 -830 840 -790
rect 1020 -830 1120 -790
<< locali >>
rect 20 200 470 210
rect 20 180 30 200
rect 110 190 470 200
rect 110 180 260 190
rect 250 170 260 180
rect 390 170 470 190
rect -430 160 0 170
rect -430 120 -50 160
rect -10 120 0 160
rect 430 150 470 170
rect 430 130 440 150
rect 460 130 470 150
rect 430 120 470 130
rect -430 110 0 120
rect -430 50 0 60
rect -430 10 -50 50
rect -10 10 0 50
rect -430 0 0 10
rect 430 40 470 50
rect 430 20 440 40
rect 460 20 470 40
rect 430 0 470 20
rect 250 -10 260 0
rect 20 -30 30 -10
rect 110 -20 260 -10
rect 390 -20 470 0
rect 110 -30 470 -20
rect 20 -40 470 -30
rect -110 -90 -100 -40
rect 170 -70 400 -60
rect 170 -90 260 -70
rect 390 -90 400 -70
rect -20 -100 120 -90
rect -20 -120 30 -100
rect 110 -120 120 -100
rect -110 -160 -100 -120
rect -430 -200 -10 -190
rect -430 -230 -40 -200
rect -430 -240 -10 -230
rect -110 -1040 -100 -270
rect 170 -350 200 -90
rect 250 -280 260 -260
rect 390 -280 400 -260
rect 250 -290 400 -280
rect 600 -290 610 200
rect 870 -130 1000 -110
rect 1020 -130 1030 -110
rect 870 -170 980 -130
rect 160 -360 210 -350
rect 160 -370 170 -360
rect 130 -390 170 -370
rect 200 -390 210 -360
rect 130 -400 210 -390
rect 310 -370 340 -290
rect 310 -400 380 -370
rect -10 -560 20 -460
rect 130 -470 160 -400
rect -10 -610 30 -560
rect -10 -630 0 -610
rect 20 -630 30 -610
rect 130 -590 160 -550
rect 350 -470 380 -400
rect 870 -450 960 -170
rect 870 -460 980 -450
rect 1090 -170 1130 -160
rect 1110 -450 1130 -170
rect 350 -580 380 -550
rect 130 -620 230 -590
rect 280 -610 300 -580
rect 330 -610 440 -580
rect -10 -640 30 -630
rect 200 -660 230 -620
rect 400 -660 440 -610
rect 200 -680 260 -660
rect 280 -680 300 -660
rect 350 -680 365 -660
rect 385 -680 440 -660
rect 240 -720 270 -710
rect 240 -800 250 -720
rect 240 -810 270 -800
rect 380 -720 410 -710
rect 400 -770 410 -720
rect 400 -780 850 -770
rect 400 -800 450 -780
rect 470 -790 850 -780
rect 470 -800 740 -790
rect 140 -820 270 -810
rect 140 -840 150 -820
rect 170 -840 270 -820
rect 140 -850 270 -840
rect 380 -830 740 -800
rect 840 -830 850 -790
rect 380 -850 850 -830
rect 240 -870 270 -850
rect 870 -870 910 -460
rect 240 -910 910 -870
rect 940 -560 980 -550
rect 940 -740 960 -560
rect 940 -900 980 -740
rect 1090 -780 1130 -450
rect 1200 -750 1210 -160
rect 1010 -790 1130 -780
rect 1010 -830 1020 -790
rect 1120 -830 1130 -790
rect 1010 -840 1130 -830
rect 150 -940 180 -930
rect 150 -1000 160 -940
rect 940 -960 1450 -900
rect 250 -1000 530 -960
rect 570 -1000 1450 -960
<< viali >>
rect 20 70 30 100
rect 30 70 110 100
rect 110 70 120 100
rect 250 70 260 100
rect 260 70 390 100
rect 390 70 400 100
rect -230 -160 -215 -40
rect -215 -160 -115 -40
rect -115 -90 -110 -40
rect -115 -120 -20 -90
rect -115 -160 -110 -120
rect 20 -230 30 -200
rect 30 -230 110 -200
rect 110 -230 120 -200
rect -230 -285 -110 -270
rect -230 -1025 -215 -285
rect -215 -1025 -115 -285
rect -115 -1025 -110 -285
rect -230 -1040 -110 -1025
rect 20 -330 30 -310
rect 30 -330 110 -310
rect 110 -330 120 -310
rect 20 -340 120 -330
rect 250 -190 260 -160
rect 260 -190 390 -160
rect 390 -190 400 -160
rect 610 185 690 200
rect 610 -275 615 185
rect 615 -275 690 185
rect 610 -290 690 -275
rect 20 -470 50 -460
rect 20 -550 30 -470
rect 30 -550 50 -470
rect 20 -560 50 -550
rect 240 -470 270 -460
rect 240 -550 270 -470
rect 240 -560 270 -550
rect 1020 -170 1050 -160
rect 1020 -450 1050 -170
rect 1020 -460 1050 -450
rect 460 -470 490 -460
rect 460 -550 480 -470
rect 480 -550 490 -470
rect 460 -560 490 -550
rect 20 -670 50 -660
rect 20 -750 30 -670
rect 30 -750 50 -670
rect 20 -760 50 -750
rect 130 -670 160 -660
rect 130 -750 150 -670
rect 150 -750 160 -670
rect 130 -760 160 -750
rect 310 -720 340 -710
rect 310 -800 340 -720
rect 310 -810 340 -800
rect 20 -870 50 -860
rect 20 -950 30 -870
rect 30 -950 50 -870
rect 20 -960 50 -950
rect 90 -870 120 -860
rect 90 -950 110 -870
rect 110 -950 120 -870
rect 1020 -560 1050 -550
rect 1020 -740 1040 -560
rect 1040 -740 1050 -560
rect 1020 -750 1050 -740
rect 1210 -175 1300 -160
rect 1210 -735 1215 -175
rect 1215 -735 1285 -175
rect 1285 -735 1300 -175
rect 1210 -750 1300 -735
rect 90 -960 120 -950
rect 150 -1020 160 -1000
rect 160 -1020 180 -1000
rect 150 -1050 180 -1020
rect 220 -940 250 -930
rect 220 -1020 240 -940
rect 240 -1020 250 -940
rect 530 -1000 570 -960
rect 220 -1030 250 -1020
<< metal1 >>
rect -400 -40 -100 300
rect 600 200 800 300
rect 600 120 610 200
rect -400 -160 -230 -40
rect -110 -80 -100 -40
rect 10 100 130 110
rect 10 70 20 100
rect 120 70 130 100
rect -110 -90 -10 -80
rect -20 -120 -10 -90
rect -110 -130 -10 -120
rect -110 -160 -100 -130
rect -400 -270 -100 -160
rect 10 -200 130 70
rect 240 100 610 120
rect 240 70 250 100
rect 400 70 610 100
rect 240 60 610 70
rect 600 -140 610 60
rect 240 -160 610 -140
rect 240 -190 250 -160
rect 400 -190 610 -160
rect 240 -200 610 -190
rect 10 -230 20 -200
rect 120 -230 130 -200
rect 10 -240 130 -230
rect -400 -1040 -230 -270
rect -110 -300 -100 -270
rect 600 -290 610 -200
rect 690 -290 800 200
rect 1200 -150 1400 300
rect -110 -310 130 -300
rect -110 -340 20 -310
rect 120 -340 130 -310
rect -110 -350 130 -340
rect -110 -650 -100 -350
rect 10 -460 500 -450
rect 10 -560 20 -460
rect 50 -560 240 -460
rect 270 -560 460 -460
rect 490 -560 500 -460
rect 10 -570 500 -560
rect -110 -660 60 -650
rect -110 -760 20 -660
rect 50 -760 60 -660
rect -110 -770 60 -760
rect 120 -660 170 -570
rect 120 -760 130 -660
rect 160 -760 170 -660
rect 120 -770 170 -760
rect 300 -710 350 -700
rect -110 -850 -100 -770
rect 300 -810 310 -710
rect 340 -810 350 -710
rect 300 -850 350 -810
rect -110 -860 60 -850
rect -110 -960 20 -860
rect 50 -960 60 -860
rect -110 -990 60 -960
rect 80 -860 350 -850
rect 80 -960 90 -860
rect 120 -900 350 -860
rect 120 -960 130 -900
rect 80 -970 130 -960
rect 210 -930 260 -920
rect -110 -1000 190 -990
rect -110 -1040 150 -1000
rect -400 -1050 150 -1040
rect 180 -1050 190 -1000
rect 210 -1030 220 -930
rect 250 -960 260 -930
rect 520 -960 580 -950
rect 250 -1000 530 -960
rect 570 -1000 580 -960
rect 250 -1030 260 -1000
rect 520 -1010 580 -1000
rect 210 -1040 260 -1030
rect -400 -1060 190 -1050
rect -400 -1100 -100 -1060
rect 600 -1100 800 -290
rect 1010 -160 1400 -150
rect 1010 -460 1020 -160
rect 1050 -460 1210 -160
rect 1010 -470 1210 -460
rect 1200 -540 1210 -470
rect 1010 -550 1210 -540
rect 1010 -750 1020 -550
rect 1050 -750 1210 -550
rect 1300 -750 1400 -160
rect 1010 -760 1400 -750
rect 1200 -1100 1400 -760
<< labels >>
rlabel metal1 -400 -1100 -100 -1080 1 VGND
port 1 n
rlabel metal1 600 -1100 800 -1080 1 VDD3v3
port 2 n
rlabel metal1 1200 -1100 1400 -1080 1 VDD1v8
port 3 n
rlabel locali 540 -800 560 -780 1 VOPAMP
rlabel locali 400 -650 420 -630 1 VOP
rlabel locali 170 190 190 210 1 VPAMP
rlabel locali 160 -30 180 -20 1 VNAMP
rlabel locali 180 -260 190 -240 1 VON
rlabel metal1 50 -70 80 -50 1 ISINK
rlabel metal1 140 -650 150 -640 1 DECISINK
rlabel locali 540 -900 570 -880 1 VONAMP
rlabel metal1 140 -890 170 -860 1 DIFFSINK
rlabel metal1 -400 280 -100 300 1 VGND
port 1 n
rlabel locali -430 110 -410 170 1 VP
port 7 n
rlabel locali -430 0 -410 60 1 VN
port 6 n
rlabel locali -430 -240 -410 -190 1 BIASN
port 5 n
rlabel locali 1430 -1000 1450 -900 1 VOUT
port 4 n
rlabel metal1 600 280 800 300 1 VDD3v3
port 2 n
rlabel metal1 1200 280 1400 300 1 VDD1v8
port 3 n
<< end >>
