magic
tech sky130A
magscale 1 2
timestamp 1635946216
<< locali >>
rect -69 17 69 33
rect -69 -17 -53 17
rect -19 -17 19 17
rect 53 -17 69 17
rect -69 -33 69 -17
<< viali >>
rect -53 -17 -19 17
rect 19 -17 53 17
<< metal1 >>
rect -65 17 65 29
rect -65 -17 -53 17
rect -19 -17 19 17
rect 53 -17 65 17
rect -65 -29 65 -17
<< end >>
