magic
tech sky130A
magscale 1 2
timestamp 1635946216
<< error_s >>
rect -2762 849 -2556 983
rect -1862 849 -1656 983
rect -962 849 -756 983
rect -62 849 144 983
rect 838 849 1044 983
rect 1738 849 1944 983
rect 2638 849 2844 983
rect 3538 849 3744 983
rect -2979 222 -2949 754
rect -2913 288 -2883 688
rect -2427 288 -2397 688
rect -2361 222 -2331 754
rect -2079 222 -2049 754
rect -2013 288 -1983 688
rect -1527 288 -1497 688
rect -1461 222 -1431 754
rect -1179 222 -1149 754
rect -1113 288 -1083 688
rect -627 288 -597 688
rect -561 222 -531 754
rect -279 222 -249 754
rect -213 288 -183 688
rect 273 288 303 688
rect 339 222 369 754
rect 621 222 651 754
rect 687 288 717 688
rect 1173 288 1203 688
rect 1239 222 1269 754
rect 1521 222 1551 754
rect 1587 288 1617 688
rect 2073 288 2103 688
rect 2139 222 2169 754
rect 2421 222 2451 754
rect 2487 288 2517 688
rect 2973 288 3003 688
rect 3039 222 3069 754
rect 3321 222 3351 754
rect 3387 288 3417 688
rect 3873 288 3903 688
rect 3939 222 3969 754
rect -2979 -518 -2949 14
rect -2913 -452 -2883 -52
rect -2427 -452 -2397 -52
rect -2361 -518 -2331 14
rect -2079 -518 -2049 14
rect -2013 -452 -1983 -52
rect -1527 -452 -1497 -52
rect -1461 -518 -1431 14
rect -1179 -518 -1149 14
rect -1113 -452 -1083 -52
rect -627 -452 -597 -52
rect -561 -518 -531 14
rect -279 -518 -249 14
rect -213 -452 -183 -52
rect 273 -452 303 -52
rect 339 -518 369 14
rect 621 -518 651 14
rect 687 -452 717 -52
rect 1173 -452 1203 -52
rect 1239 -518 1269 14
rect 1521 -518 1551 14
rect 1587 -452 1617 -52
rect 2073 -452 2103 -52
rect 2139 -518 2169 14
rect 2421 -518 2451 14
rect 2487 -452 2517 -52
rect 2973 -452 3003 -52
rect 3039 -518 3069 14
rect 3321 -518 3351 14
rect 3387 -452 3417 -52
rect 3873 -452 3903 -52
rect 3939 -518 3969 14
rect -2765 -756 -2559 -622
rect -1865 -756 -1659 -622
rect -965 -756 -759 -622
rect -65 -756 141 -622
rect 835 -756 1041 -622
rect 1735 -756 1941 -622
rect 2635 -756 2841 -622
rect 3535 -756 3741 -622
<< metal1 >>
rect -3371 1130 3393 1313
rect -2403 -1097 4030 -911
<< metal2 >>
rect -2759 68 3734 168
use contact$4  contact$4_0
array 0 7 900 0 0 0
timestamp 1635946216
transform 1 0 -2645 0 1 118
box -64 -32 64 32
use m2_pfet_w2_l2  m2_pfet_w2_l2_0
array 0 7 900 0 0 0
timestamp 1635946216
transform 1 0 -2655 0 1 -252
box -385 -659 385 1382
<< end >>
