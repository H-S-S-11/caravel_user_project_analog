magic
tech sky130A
magscale 1 2
timestamp 1632242116
<< nwell >>
rect -545 -447 545 447
<< mvpmos >>
rect -287 -150 -187 150
rect -129 -150 -29 150
rect 29 -150 129 150
rect 187 -150 287 150
<< mvpdiff >>
rect -345 138 -287 150
rect -345 -138 -333 138
rect -299 -138 -287 138
rect -345 -150 -287 -138
rect -187 138 -129 150
rect -187 -138 -175 138
rect -141 -138 -129 138
rect -187 -150 -129 -138
rect -29 138 29 150
rect -29 -138 -17 138
rect 17 -138 29 138
rect -29 -150 29 -138
rect 129 138 187 150
rect 129 -138 141 138
rect 175 -138 187 138
rect 129 -150 187 -138
rect 287 138 345 150
rect 287 -138 299 138
rect 333 -138 345 138
rect 287 -150 345 -138
<< mvpdiffc >>
rect -333 -138 -299 138
rect -175 -138 -141 138
rect -17 -138 17 138
rect 141 -138 175 138
rect 299 -138 333 138
<< mvnsubdiff >>
rect -479 369 479 381
rect -479 335 -371 369
rect 371 335 479 369
rect -479 323 479 335
rect -479 273 -421 323
rect -479 -273 -467 273
rect -433 -273 -421 273
rect 421 273 479 323
rect -479 -323 -421 -273
rect 421 -273 433 273
rect 467 -273 479 273
rect 421 -323 479 -273
rect -479 -335 479 -323
rect -479 -369 -371 -335
rect 371 -369 479 -335
rect -479 -381 479 -369
<< mvnsubdiffcont >>
rect -371 335 371 369
rect -467 -273 -433 273
rect 433 -273 467 273
rect -371 -369 371 -335
<< poly >>
rect -287 231 -187 247
rect -287 197 -271 231
rect -203 197 -187 231
rect -287 150 -187 197
rect -129 231 -29 247
rect -129 197 -113 231
rect -45 197 -29 231
rect -129 150 -29 197
rect 29 231 129 247
rect 29 197 45 231
rect 113 197 129 231
rect 29 150 129 197
rect 187 231 287 247
rect 187 197 203 231
rect 271 197 287 231
rect 187 150 287 197
rect -287 -197 -187 -150
rect -287 -231 -271 -197
rect -203 -231 -187 -197
rect -287 -247 -187 -231
rect -129 -197 -29 -150
rect -129 -231 -113 -197
rect -45 -231 -29 -197
rect -129 -247 -29 -231
rect 29 -197 129 -150
rect 29 -231 45 -197
rect 113 -231 129 -197
rect 29 -247 129 -231
rect 187 -197 287 -150
rect 187 -231 203 -197
rect 271 -231 287 -197
rect 187 -247 287 -231
<< polycont >>
rect -271 197 -203 231
rect -113 197 -45 231
rect 45 197 113 231
rect 203 197 271 231
rect -271 -231 -203 -197
rect -113 -231 -45 -197
rect 45 -231 113 -197
rect 203 -231 271 -197
<< locali >>
rect -467 335 -371 369
rect 371 335 467 369
rect -467 273 -433 335
rect 433 273 467 335
rect -287 197 -271 231
rect -203 197 -187 231
rect -129 197 -113 231
rect -45 197 -29 231
rect 29 197 45 231
rect 113 197 129 231
rect 187 197 203 231
rect 271 197 287 231
rect -333 138 -299 154
rect -333 -154 -299 -138
rect -175 138 -141 154
rect -175 -154 -141 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 141 138 175 154
rect 141 -154 175 -138
rect 299 138 333 154
rect 299 -154 333 -138
rect -287 -231 -271 -197
rect -203 -231 -187 -197
rect -129 -231 -113 -197
rect -45 -231 -29 -197
rect 29 -231 45 -197
rect 113 -231 129 -197
rect 187 -231 203 -197
rect 271 -231 287 -197
rect -467 -335 -433 -273
rect 433 -335 467 -273
rect -467 -369 -371 -335
rect 371 -369 467 -335
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string FIXED_BBOX -450 -352 450 352
string parameters w 1.5 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
