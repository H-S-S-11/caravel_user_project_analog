magic
tech sky130A
magscale 1 2
timestamp 1635946216
<< error_s >>
rect -2830 2113 -2604 2149
rect -2830 2031 -2794 2113
rect -2640 2031 -2604 2113
rect -2830 1995 -2604 2031
rect -2746 1832 -2744 1866
rect -2710 1832 -2706 1866
rect -2872 1728 -2838 1730
rect -2614 1728 -2580 1730
rect -2872 1712 -2838 1714
rect -2614 1712 -2580 1714
rect -2872 1674 -2838 1676
rect -2614 1674 -2580 1676
rect -2872 1660 -2838 1662
rect -2614 1660 -2580 1662
rect -2872 1640 -2838 1642
rect -2614 1640 -2580 1642
rect -2872 1602 -2838 1604
rect -2614 1602 -2580 1604
rect -2872 1592 -2838 1594
rect -2614 1592 -2580 1594
rect -2872 1568 -2838 1570
rect -2614 1568 -2580 1570
rect -2872 1530 -2838 1532
rect -2614 1530 -2580 1532
rect -2872 1524 -2838 1526
rect -2614 1524 -2580 1526
rect -2872 1496 -2838 1498
rect -2614 1496 -2580 1498
rect -2872 1456 -2838 1460
rect -2614 1456 -2580 1460
rect -2872 1424 -2838 1426
rect -2614 1424 -2580 1426
rect -2872 1386 -2838 1390
rect -2614 1386 -2580 1390
rect -2872 1352 -2838 1354
rect -2614 1352 -2580 1354
rect -2872 1320 -2838 1322
rect -2614 1320 -2580 1322
rect -2872 1314 -2838 1316
rect -2614 1314 -2580 1316
rect -2872 1280 -2838 1282
rect -2614 1280 -2580 1282
rect -2872 1252 -2838 1254
rect -2614 1252 -2580 1254
rect -2872 1242 -2838 1244
rect -2614 1242 -2580 1244
rect -2872 1208 -2838 1210
rect -2614 1208 -2580 1210
rect -2872 1184 -2838 1186
rect -2614 1184 -2580 1186
rect -2872 1170 -2838 1172
rect -2614 1170 -2580 1172
rect -2872 1136 -2838 1138
rect -2614 1136 -2580 1138
rect -2872 1116 -2838 1118
rect -2614 1116 -2580 1118
rect -2872 1098 -2838 1100
rect -2614 1098 -2580 1100
rect -2872 1064 -2838 1066
rect -2614 1064 -2580 1066
rect -2872 1048 -2838 1050
rect -2614 1048 -2580 1050
rect -2872 1026 -2838 1028
rect -2614 1026 -2580 1028
rect -2872 992 -2838 994
rect -2614 992 -2580 994
rect -2872 980 -2838 982
rect -2614 980 -2580 982
rect -2872 954 -2838 956
rect -2614 954 -2580 956
rect -2872 920 -2838 922
rect -2614 920 -2580 922
rect -2872 912 -2838 914
rect -2614 912 -2580 914
rect -2872 882 -2838 884
rect -2614 882 -2580 884
rect -2872 848 -2838 850
rect -2614 848 -2580 850
rect -2872 844 -2838 846
rect -2614 844 -2580 846
rect -2872 810 -2838 812
rect -2614 810 -2580 812
rect -2872 776 -2838 778
rect -2614 776 -2580 778
rect -2872 738 -2838 740
rect -2614 738 -2580 740
rect -2872 708 -2838 710
rect -2614 708 -2580 710
rect -2872 704 -2838 706
rect -2614 704 -2580 706
rect -2872 666 -2838 668
rect -2614 666 -2580 668
rect -2872 640 -2838 642
rect -2614 640 -2580 642
rect -2872 632 -2838 634
rect -2614 632 -2580 634
rect -2872 594 -2838 596
rect -2614 594 -2580 596
rect -2872 572 -2838 574
rect -2614 572 -2580 574
rect -2872 560 -2838 562
rect -2614 560 -2580 562
rect -2872 522 -2838 524
rect -2614 522 -2580 524
rect -2872 504 -2838 506
rect -2614 504 -2580 506
rect -2872 488 -2838 490
rect -2614 488 -2580 490
rect -2872 450 -2838 452
rect -2614 450 -2580 452
rect -2872 436 -2838 438
rect -2614 436 -2580 438
rect -2872 416 -2838 418
rect -2614 416 -2580 418
rect -2872 378 -2838 380
rect -2614 378 -2580 380
rect -2872 368 -2838 370
rect -2614 368 -2580 370
rect -2872 344 -2838 346
rect -2614 344 -2580 346
rect -2872 306 -2838 308
rect -2614 306 -2580 308
rect -2872 300 -2838 302
rect -2614 300 -2580 302
rect -2872 272 -2838 274
rect -2614 272 -2580 274
rect -2872 232 -2838 236
rect -2614 232 -2580 236
rect -2872 200 -2838 202
rect -2614 200 -2580 202
rect -2872 162 -2838 166
rect -2614 162 -2580 166
rect -2872 128 -2838 130
rect -2614 128 -2580 130
rect -2872 96 -2838 98
rect -2614 96 -2580 98
rect -2872 90 -2838 92
rect -2614 90 -2580 92
rect -2872 56 -2838 58
rect -2614 56 -2580 58
rect -2872 28 -2838 30
rect -2614 28 -2580 30
rect -2872 18 -2838 20
rect -2614 18 -2580 20
rect -2872 -16 -2838 -14
rect -2614 -16 -2580 -14
rect -2872 -40 -2838 -38
rect -2614 -40 -2580 -38
rect -2872 -54 -2838 -52
rect -2614 -54 -2580 -52
rect -2872 -88 -2838 -86
rect -2614 -88 -2580 -86
rect -2872 -108 -2838 -106
rect -2614 -108 -2580 -106
rect -2872 -126 -2838 -124
rect -2614 -126 -2580 -124
rect -2746 -278 -2744 -244
rect -2710 -278 -2706 -244
<< pdiff >>
rect -2794 2031 -2640 2113
<< metal1 >>
rect -3014 -206 -2878 2344
rect -2822 -479 -2630 -284
rect -2574 -756 -2438 1794
use contact$4  contact$4_0
timestamp 1635946216
transform 1 0 -2725 0 1 -379
box -64 -32 64 32
use contact$2  contact$2_0
timestamp 1635946216
transform 1 0 -2717 0 1 2072
box -103 -67 103 67
use sky130_fd_pr__nfet_g5v0d10v5_9A4VCP  sky130_fd_pr__nfet_g5v0d10v5_9A4VCP_0
timestamp 1635946216
transform 1 0 -2726 0 1 794
box -184 -1088 184 1088
<< end >>
