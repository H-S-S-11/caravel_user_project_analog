magic
tech sky130A
magscale 1 2
timestamp 1635946216
<< error_s >>
rect -2458 2212 -2232 2248
rect -2458 2130 -2422 2212
rect -2268 2130 -2232 2212
rect -2458 2094 -2232 2130
rect -1758 2212 -1532 2248
rect -1758 2130 -1722 2212
rect -1568 2130 -1532 2212
rect -1758 2094 -1532 2130
rect -1058 2212 -832 2248
rect -1058 2130 -1022 2212
rect -868 2130 -832 2212
rect -1058 2094 -832 2130
rect -358 2212 -132 2248
rect -358 2130 -322 2212
rect -168 2130 -132 2212
rect -358 2094 -132 2130
rect 342 2212 568 2248
rect 342 2130 378 2212
rect 532 2130 568 2212
rect 342 2094 568 2130
rect 1042 2212 1268 2248
rect 1042 2130 1078 2212
rect 1232 2130 1268 2212
rect 1042 2094 1268 2130
rect 1742 2212 1968 2248
rect 1742 2130 1778 2212
rect 1932 2130 1968 2212
rect 1742 2094 1968 2130
rect 2442 2212 2668 2248
rect 2442 2130 2478 2212
rect 2632 2130 2668 2212
rect 2442 2094 2668 2130
rect 3142 2212 3368 2248
rect 3142 2130 3178 2212
rect 3332 2130 3368 2212
rect 3142 2094 3368 2130
rect 3842 2212 4068 2248
rect 3842 2130 3878 2212
rect 4032 2130 4068 2212
rect 3842 2094 4068 2130
rect -2374 1931 -2372 1965
rect -2338 1931 -2334 1965
rect -1674 1931 -1672 1965
rect -1638 1931 -1634 1965
rect -974 1931 -972 1965
rect -938 1931 -934 1965
rect -274 1931 -272 1965
rect -238 1931 -234 1965
rect 426 1931 428 1965
rect 462 1931 466 1965
rect 1126 1931 1128 1965
rect 1162 1931 1166 1965
rect 1826 1931 1828 1965
rect 1862 1931 1866 1965
rect 2526 1931 2528 1965
rect 2562 1931 2566 1965
rect 3226 1931 3228 1965
rect 3262 1931 3266 1965
rect 3926 1931 3928 1965
rect 3962 1931 3966 1965
rect -2500 1827 -2466 1829
rect -2242 1827 -2208 1829
rect -1800 1827 -1766 1829
rect -1542 1827 -1508 1829
rect -1100 1827 -1066 1829
rect -842 1827 -808 1829
rect -400 1827 -366 1829
rect -142 1827 -108 1829
rect 300 1827 334 1829
rect 558 1827 592 1829
rect 1000 1827 1034 1829
rect 1258 1827 1292 1829
rect 1700 1827 1734 1829
rect 1958 1827 1992 1829
rect 2400 1827 2434 1829
rect 2658 1827 2692 1829
rect 3100 1827 3134 1829
rect 3358 1827 3392 1829
rect 3800 1827 3834 1829
rect 4058 1827 4092 1829
rect -2500 1811 -2466 1813
rect -2242 1811 -2208 1813
rect -1800 1811 -1766 1813
rect -1542 1811 -1508 1813
rect -1100 1811 -1066 1813
rect -842 1811 -808 1813
rect -400 1811 -366 1813
rect -142 1811 -108 1813
rect 300 1811 334 1813
rect 558 1811 592 1813
rect 1000 1811 1034 1813
rect 1258 1811 1292 1813
rect 1700 1811 1734 1813
rect 1958 1811 1992 1813
rect 2400 1811 2434 1813
rect 2658 1811 2692 1813
rect 3100 1811 3134 1813
rect 3358 1811 3392 1813
rect 3800 1811 3834 1813
rect 4058 1811 4092 1813
rect -2500 1773 -2466 1775
rect -2242 1773 -2208 1775
rect -1800 1773 -1766 1775
rect -1542 1773 -1508 1775
rect -1100 1773 -1066 1775
rect -842 1773 -808 1775
rect -400 1773 -366 1775
rect -142 1773 -108 1775
rect 300 1773 334 1775
rect 558 1773 592 1775
rect 1000 1773 1034 1775
rect 1258 1773 1292 1775
rect 1700 1773 1734 1775
rect 1958 1773 1992 1775
rect 2400 1773 2434 1775
rect 2658 1773 2692 1775
rect 3100 1773 3134 1775
rect 3358 1773 3392 1775
rect 3800 1773 3834 1775
rect 4058 1773 4092 1775
rect -2500 1759 -2466 1761
rect -2242 1759 -2208 1761
rect -1800 1759 -1766 1761
rect -1542 1759 -1508 1761
rect -1100 1759 -1066 1761
rect -842 1759 -808 1761
rect -400 1759 -366 1761
rect -142 1759 -108 1761
rect 300 1759 334 1761
rect 558 1759 592 1761
rect 1000 1759 1034 1761
rect 1258 1759 1292 1761
rect 1700 1759 1734 1761
rect 1958 1759 1992 1761
rect 2400 1759 2434 1761
rect 2658 1759 2692 1761
rect 3100 1759 3134 1761
rect 3358 1759 3392 1761
rect 3800 1759 3834 1761
rect 4058 1759 4092 1761
rect -2500 1739 -2466 1741
rect -2242 1739 -2208 1741
rect -1800 1739 -1766 1741
rect -1542 1739 -1508 1741
rect -1100 1739 -1066 1741
rect -842 1739 -808 1741
rect -400 1739 -366 1741
rect -142 1739 -108 1741
rect 300 1739 334 1741
rect 558 1739 592 1741
rect 1000 1739 1034 1741
rect 1258 1739 1292 1741
rect 1700 1739 1734 1741
rect 1958 1739 1992 1741
rect 2400 1739 2434 1741
rect 2658 1739 2692 1741
rect 3100 1739 3134 1741
rect 3358 1739 3392 1741
rect 3800 1739 3834 1741
rect 4058 1739 4092 1741
rect -2500 1701 -2466 1703
rect -2242 1701 -2208 1703
rect -1800 1701 -1766 1703
rect -1542 1701 -1508 1703
rect -1100 1701 -1066 1703
rect -842 1701 -808 1703
rect -400 1701 -366 1703
rect -142 1701 -108 1703
rect 300 1701 334 1703
rect 558 1701 592 1703
rect 1000 1701 1034 1703
rect 1258 1701 1292 1703
rect 1700 1701 1734 1703
rect 1958 1701 1992 1703
rect 2400 1701 2434 1703
rect 2658 1701 2692 1703
rect 3100 1701 3134 1703
rect 3358 1701 3392 1703
rect 3800 1701 3834 1703
rect 4058 1701 4092 1703
rect -2500 1691 -2466 1693
rect -2242 1691 -2208 1693
rect -1800 1691 -1766 1693
rect -1542 1691 -1508 1693
rect -1100 1691 -1066 1693
rect -842 1691 -808 1693
rect -400 1691 -366 1693
rect -142 1691 -108 1693
rect 300 1691 334 1693
rect 558 1691 592 1693
rect 1000 1691 1034 1693
rect 1258 1691 1292 1693
rect 1700 1691 1734 1693
rect 1958 1691 1992 1693
rect 2400 1691 2434 1693
rect 2658 1691 2692 1693
rect 3100 1691 3134 1693
rect 3358 1691 3392 1693
rect 3800 1691 3834 1693
rect 4058 1691 4092 1693
rect -2500 1667 -2466 1669
rect -2242 1667 -2208 1669
rect -1800 1667 -1766 1669
rect -1542 1667 -1508 1669
rect -1100 1667 -1066 1669
rect -842 1667 -808 1669
rect -400 1667 -366 1669
rect -142 1667 -108 1669
rect 300 1667 334 1669
rect 558 1667 592 1669
rect 1000 1667 1034 1669
rect 1258 1667 1292 1669
rect 1700 1667 1734 1669
rect 1958 1667 1992 1669
rect 2400 1667 2434 1669
rect 2658 1667 2692 1669
rect 3100 1667 3134 1669
rect 3358 1667 3392 1669
rect 3800 1667 3834 1669
rect 4058 1667 4092 1669
rect -2500 1629 -2466 1631
rect -2242 1629 -2208 1631
rect -1800 1629 -1766 1631
rect -1542 1629 -1508 1631
rect -1100 1629 -1066 1631
rect -842 1629 -808 1631
rect -400 1629 -366 1631
rect -142 1629 -108 1631
rect 300 1629 334 1631
rect 558 1629 592 1631
rect 1000 1629 1034 1631
rect 1258 1629 1292 1631
rect 1700 1629 1734 1631
rect 1958 1629 1992 1631
rect 2400 1629 2434 1631
rect 2658 1629 2692 1631
rect 3100 1629 3134 1631
rect 3358 1629 3392 1631
rect 3800 1629 3834 1631
rect 4058 1629 4092 1631
rect -2500 1623 -2466 1625
rect -2242 1623 -2208 1625
rect -1800 1623 -1766 1625
rect -1542 1623 -1508 1625
rect -1100 1623 -1066 1625
rect -842 1623 -808 1625
rect -400 1623 -366 1625
rect -142 1623 -108 1625
rect 300 1623 334 1625
rect 558 1623 592 1625
rect 1000 1623 1034 1625
rect 1258 1623 1292 1625
rect 1700 1623 1734 1625
rect 1958 1623 1992 1625
rect 2400 1623 2434 1625
rect 2658 1623 2692 1625
rect 3100 1623 3134 1625
rect 3358 1623 3392 1625
rect 3800 1623 3834 1625
rect 4058 1623 4092 1625
rect -2500 1595 -2466 1597
rect -2242 1595 -2208 1597
rect -1800 1595 -1766 1597
rect -1542 1595 -1508 1597
rect -1100 1595 -1066 1597
rect -842 1595 -808 1597
rect -400 1595 -366 1597
rect -142 1595 -108 1597
rect 300 1595 334 1597
rect 558 1595 592 1597
rect 1000 1595 1034 1597
rect 1258 1595 1292 1597
rect 1700 1595 1734 1597
rect 1958 1595 1992 1597
rect 2400 1595 2434 1597
rect 2658 1595 2692 1597
rect 3100 1595 3134 1597
rect 3358 1595 3392 1597
rect 3800 1595 3834 1597
rect 4058 1595 4092 1597
rect -2500 1555 -2466 1559
rect -2242 1555 -2208 1559
rect -1800 1555 -1766 1559
rect -1542 1555 -1508 1559
rect -1100 1555 -1066 1559
rect -842 1555 -808 1559
rect -400 1555 -366 1559
rect -142 1555 -108 1559
rect 300 1555 334 1559
rect 558 1555 592 1559
rect 1000 1555 1034 1559
rect 1258 1555 1292 1559
rect 1700 1555 1734 1559
rect 1958 1555 1992 1559
rect 2400 1555 2434 1559
rect 2658 1555 2692 1559
rect 3100 1555 3134 1559
rect 3358 1555 3392 1559
rect 3800 1555 3834 1559
rect 4058 1555 4092 1559
rect -2500 1523 -2466 1525
rect -2242 1523 -2208 1525
rect -1800 1523 -1766 1525
rect -1542 1523 -1508 1525
rect -1100 1523 -1066 1525
rect -842 1523 -808 1525
rect -400 1523 -366 1525
rect -142 1523 -108 1525
rect 300 1523 334 1525
rect 558 1523 592 1525
rect 1000 1523 1034 1525
rect 1258 1523 1292 1525
rect 1700 1523 1734 1525
rect 1958 1523 1992 1525
rect 2400 1523 2434 1525
rect 2658 1523 2692 1525
rect 3100 1523 3134 1525
rect 3358 1523 3392 1525
rect 3800 1523 3834 1525
rect 4058 1523 4092 1525
rect -2500 1485 -2466 1489
rect -2242 1485 -2208 1489
rect -1800 1485 -1766 1489
rect -1542 1485 -1508 1489
rect -1100 1485 -1066 1489
rect -842 1485 -808 1489
rect -400 1485 -366 1489
rect -142 1485 -108 1489
rect 300 1485 334 1489
rect 558 1485 592 1489
rect 1000 1485 1034 1489
rect 1258 1485 1292 1489
rect 1700 1485 1734 1489
rect 1958 1485 1992 1489
rect 2400 1485 2434 1489
rect 2658 1485 2692 1489
rect 3100 1485 3134 1489
rect 3358 1485 3392 1489
rect 3800 1485 3834 1489
rect 4058 1485 4092 1489
rect -2500 1451 -2466 1453
rect -2242 1451 -2208 1453
rect -1800 1451 -1766 1453
rect -1542 1451 -1508 1453
rect -1100 1451 -1066 1453
rect -842 1451 -808 1453
rect -400 1451 -366 1453
rect -142 1451 -108 1453
rect 300 1451 334 1453
rect 558 1451 592 1453
rect 1000 1451 1034 1453
rect 1258 1451 1292 1453
rect 1700 1451 1734 1453
rect 1958 1451 1992 1453
rect 2400 1451 2434 1453
rect 2658 1451 2692 1453
rect 3100 1451 3134 1453
rect 3358 1451 3392 1453
rect 3800 1451 3834 1453
rect 4058 1451 4092 1453
rect -2500 1419 -2466 1421
rect -2242 1419 -2208 1421
rect -1800 1419 -1766 1421
rect -1542 1419 -1508 1421
rect -1100 1419 -1066 1421
rect -842 1419 -808 1421
rect -400 1419 -366 1421
rect -142 1419 -108 1421
rect 300 1419 334 1421
rect 558 1419 592 1421
rect 1000 1419 1034 1421
rect 1258 1419 1292 1421
rect 1700 1419 1734 1421
rect 1958 1419 1992 1421
rect 2400 1419 2434 1421
rect 2658 1419 2692 1421
rect 3100 1419 3134 1421
rect 3358 1419 3392 1421
rect 3800 1419 3834 1421
rect 4058 1419 4092 1421
rect -2500 1413 -2466 1415
rect -2242 1413 -2208 1415
rect -1800 1413 -1766 1415
rect -1542 1413 -1508 1415
rect -1100 1413 -1066 1415
rect -842 1413 -808 1415
rect -400 1413 -366 1415
rect -142 1413 -108 1415
rect 300 1413 334 1415
rect 558 1413 592 1415
rect 1000 1413 1034 1415
rect 1258 1413 1292 1415
rect 1700 1413 1734 1415
rect 1958 1413 1992 1415
rect 2400 1413 2434 1415
rect 2658 1413 2692 1415
rect 3100 1413 3134 1415
rect 3358 1413 3392 1415
rect 3800 1413 3834 1415
rect 4058 1413 4092 1415
rect -2500 1379 -2466 1381
rect -2242 1379 -2208 1381
rect -1800 1379 -1766 1381
rect -1542 1379 -1508 1381
rect -1100 1379 -1066 1381
rect -842 1379 -808 1381
rect -400 1379 -366 1381
rect -142 1379 -108 1381
rect 300 1379 334 1381
rect 558 1379 592 1381
rect 1000 1379 1034 1381
rect 1258 1379 1292 1381
rect 1700 1379 1734 1381
rect 1958 1379 1992 1381
rect 2400 1379 2434 1381
rect 2658 1379 2692 1381
rect 3100 1379 3134 1381
rect 3358 1379 3392 1381
rect 3800 1379 3834 1381
rect 4058 1379 4092 1381
rect -2500 1351 -2466 1353
rect -2242 1351 -2208 1353
rect -1800 1351 -1766 1353
rect -1542 1351 -1508 1353
rect -1100 1351 -1066 1353
rect -842 1351 -808 1353
rect -400 1351 -366 1353
rect -142 1351 -108 1353
rect 300 1351 334 1353
rect 558 1351 592 1353
rect 1000 1351 1034 1353
rect 1258 1351 1292 1353
rect 1700 1351 1734 1353
rect 1958 1351 1992 1353
rect 2400 1351 2434 1353
rect 2658 1351 2692 1353
rect 3100 1351 3134 1353
rect 3358 1351 3392 1353
rect 3800 1351 3834 1353
rect 4058 1351 4092 1353
rect -2500 1341 -2466 1343
rect -2242 1341 -2208 1343
rect -1800 1341 -1766 1343
rect -1542 1341 -1508 1343
rect -1100 1341 -1066 1343
rect -842 1341 -808 1343
rect -400 1341 -366 1343
rect -142 1341 -108 1343
rect 300 1341 334 1343
rect 558 1341 592 1343
rect 1000 1341 1034 1343
rect 1258 1341 1292 1343
rect 1700 1341 1734 1343
rect 1958 1341 1992 1343
rect 2400 1341 2434 1343
rect 2658 1341 2692 1343
rect 3100 1341 3134 1343
rect 3358 1341 3392 1343
rect 3800 1341 3834 1343
rect 4058 1341 4092 1343
rect -2500 1307 -2466 1309
rect -2242 1307 -2208 1309
rect -1800 1307 -1766 1309
rect -1542 1307 -1508 1309
rect -1100 1307 -1066 1309
rect -842 1307 -808 1309
rect -400 1307 -366 1309
rect -142 1307 -108 1309
rect 300 1307 334 1309
rect 558 1307 592 1309
rect 1000 1307 1034 1309
rect 1258 1307 1292 1309
rect 1700 1307 1734 1309
rect 1958 1307 1992 1309
rect 2400 1307 2434 1309
rect 2658 1307 2692 1309
rect 3100 1307 3134 1309
rect 3358 1307 3392 1309
rect 3800 1307 3834 1309
rect 4058 1307 4092 1309
rect -2500 1283 -2466 1285
rect -2242 1283 -2208 1285
rect -1800 1283 -1766 1285
rect -1542 1283 -1508 1285
rect -1100 1283 -1066 1285
rect -842 1283 -808 1285
rect -400 1283 -366 1285
rect -142 1283 -108 1285
rect 300 1283 334 1285
rect 558 1283 592 1285
rect 1000 1283 1034 1285
rect 1258 1283 1292 1285
rect 1700 1283 1734 1285
rect 1958 1283 1992 1285
rect 2400 1283 2434 1285
rect 2658 1283 2692 1285
rect 3100 1283 3134 1285
rect 3358 1283 3392 1285
rect 3800 1283 3834 1285
rect 4058 1283 4092 1285
rect -2500 1269 -2466 1271
rect -2242 1269 -2208 1271
rect -1800 1269 -1766 1271
rect -1542 1269 -1508 1271
rect -1100 1269 -1066 1271
rect -842 1269 -808 1271
rect -400 1269 -366 1271
rect -142 1269 -108 1271
rect 300 1269 334 1271
rect 558 1269 592 1271
rect 1000 1269 1034 1271
rect 1258 1269 1292 1271
rect 1700 1269 1734 1271
rect 1958 1269 1992 1271
rect 2400 1269 2434 1271
rect 2658 1269 2692 1271
rect 3100 1269 3134 1271
rect 3358 1269 3392 1271
rect 3800 1269 3834 1271
rect 4058 1269 4092 1271
rect -2500 1235 -2466 1237
rect -2242 1235 -2208 1237
rect -1800 1235 -1766 1237
rect -1542 1235 -1508 1237
rect -1100 1235 -1066 1237
rect -842 1235 -808 1237
rect -400 1235 -366 1237
rect -142 1235 -108 1237
rect 300 1235 334 1237
rect 558 1235 592 1237
rect 1000 1235 1034 1237
rect 1258 1235 1292 1237
rect 1700 1235 1734 1237
rect 1958 1235 1992 1237
rect 2400 1235 2434 1237
rect 2658 1235 2692 1237
rect 3100 1235 3134 1237
rect 3358 1235 3392 1237
rect 3800 1235 3834 1237
rect 4058 1235 4092 1237
rect -2500 1215 -2466 1217
rect -2242 1215 -2208 1217
rect -1800 1215 -1766 1217
rect -1542 1215 -1508 1217
rect -1100 1215 -1066 1217
rect -842 1215 -808 1217
rect -400 1215 -366 1217
rect -142 1215 -108 1217
rect 300 1215 334 1217
rect 558 1215 592 1217
rect 1000 1215 1034 1217
rect 1258 1215 1292 1217
rect 1700 1215 1734 1217
rect 1958 1215 1992 1217
rect 2400 1215 2434 1217
rect 2658 1215 2692 1217
rect 3100 1215 3134 1217
rect 3358 1215 3392 1217
rect 3800 1215 3834 1217
rect 4058 1215 4092 1217
rect -2500 1197 -2466 1199
rect -2242 1197 -2208 1199
rect -1800 1197 -1766 1199
rect -1542 1197 -1508 1199
rect -1100 1197 -1066 1199
rect -842 1197 -808 1199
rect -400 1197 -366 1199
rect -142 1197 -108 1199
rect 300 1197 334 1199
rect 558 1197 592 1199
rect 1000 1197 1034 1199
rect 1258 1197 1292 1199
rect 1700 1197 1734 1199
rect 1958 1197 1992 1199
rect 2400 1197 2434 1199
rect 2658 1197 2692 1199
rect 3100 1197 3134 1199
rect 3358 1197 3392 1199
rect 3800 1197 3834 1199
rect 4058 1197 4092 1199
rect -2500 1163 -2466 1165
rect -2242 1163 -2208 1165
rect -1800 1163 -1766 1165
rect -1542 1163 -1508 1165
rect -1100 1163 -1066 1165
rect -842 1163 -808 1165
rect -400 1163 -366 1165
rect -142 1163 -108 1165
rect 300 1163 334 1165
rect 558 1163 592 1165
rect 1000 1163 1034 1165
rect 1258 1163 1292 1165
rect 1700 1163 1734 1165
rect 1958 1163 1992 1165
rect 2400 1163 2434 1165
rect 2658 1163 2692 1165
rect 3100 1163 3134 1165
rect 3358 1163 3392 1165
rect 3800 1163 3834 1165
rect 4058 1163 4092 1165
rect -2500 1147 -2466 1149
rect -2242 1147 -2208 1149
rect -1800 1147 -1766 1149
rect -1542 1147 -1508 1149
rect -1100 1147 -1066 1149
rect -842 1147 -808 1149
rect -400 1147 -366 1149
rect -142 1147 -108 1149
rect 300 1147 334 1149
rect 558 1147 592 1149
rect 1000 1147 1034 1149
rect 1258 1147 1292 1149
rect 1700 1147 1734 1149
rect 1958 1147 1992 1149
rect 2400 1147 2434 1149
rect 2658 1147 2692 1149
rect 3100 1147 3134 1149
rect 3358 1147 3392 1149
rect 3800 1147 3834 1149
rect 4058 1147 4092 1149
rect -2500 1125 -2466 1127
rect -2242 1125 -2208 1127
rect -1800 1125 -1766 1127
rect -1542 1125 -1508 1127
rect -1100 1125 -1066 1127
rect -842 1125 -808 1127
rect -400 1125 -366 1127
rect -142 1125 -108 1127
rect 300 1125 334 1127
rect 558 1125 592 1127
rect 1000 1125 1034 1127
rect 1258 1125 1292 1127
rect 1700 1125 1734 1127
rect 1958 1125 1992 1127
rect 2400 1125 2434 1127
rect 2658 1125 2692 1127
rect 3100 1125 3134 1127
rect 3358 1125 3392 1127
rect 3800 1125 3834 1127
rect 4058 1125 4092 1127
rect -2500 1091 -2466 1093
rect -2242 1091 -2208 1093
rect -1800 1091 -1766 1093
rect -1542 1091 -1508 1093
rect -1100 1091 -1066 1093
rect -842 1091 -808 1093
rect -400 1091 -366 1093
rect -142 1091 -108 1093
rect 300 1091 334 1093
rect 558 1091 592 1093
rect 1000 1091 1034 1093
rect 1258 1091 1292 1093
rect 1700 1091 1734 1093
rect 1958 1091 1992 1093
rect 2400 1091 2434 1093
rect 2658 1091 2692 1093
rect 3100 1091 3134 1093
rect 3358 1091 3392 1093
rect 3800 1091 3834 1093
rect 4058 1091 4092 1093
rect -2500 1079 -2466 1081
rect -2242 1079 -2208 1081
rect -1800 1079 -1766 1081
rect -1542 1079 -1508 1081
rect -1100 1079 -1066 1081
rect -842 1079 -808 1081
rect -400 1079 -366 1081
rect -142 1079 -108 1081
rect 300 1079 334 1081
rect 558 1079 592 1081
rect 1000 1079 1034 1081
rect 1258 1079 1292 1081
rect 1700 1079 1734 1081
rect 1958 1079 1992 1081
rect 2400 1079 2434 1081
rect 2658 1079 2692 1081
rect 3100 1079 3134 1081
rect 3358 1079 3392 1081
rect 3800 1079 3834 1081
rect 4058 1079 4092 1081
rect -2500 1053 -2466 1055
rect -2242 1053 -2208 1055
rect -1800 1053 -1766 1055
rect -1542 1053 -1508 1055
rect -1100 1053 -1066 1055
rect -842 1053 -808 1055
rect -400 1053 -366 1055
rect -142 1053 -108 1055
rect 300 1053 334 1055
rect 558 1053 592 1055
rect 1000 1053 1034 1055
rect 1258 1053 1292 1055
rect 1700 1053 1734 1055
rect 1958 1053 1992 1055
rect 2400 1053 2434 1055
rect 2658 1053 2692 1055
rect 3100 1053 3134 1055
rect 3358 1053 3392 1055
rect 3800 1053 3834 1055
rect 4058 1053 4092 1055
rect -2500 1019 -2466 1021
rect -2242 1019 -2208 1021
rect -1800 1019 -1766 1021
rect -1542 1019 -1508 1021
rect -1100 1019 -1066 1021
rect -842 1019 -808 1021
rect -400 1019 -366 1021
rect -142 1019 -108 1021
rect 300 1019 334 1021
rect 558 1019 592 1021
rect 1000 1019 1034 1021
rect 1258 1019 1292 1021
rect 1700 1019 1734 1021
rect 1958 1019 1992 1021
rect 2400 1019 2434 1021
rect 2658 1019 2692 1021
rect 3100 1019 3134 1021
rect 3358 1019 3392 1021
rect 3800 1019 3834 1021
rect 4058 1019 4092 1021
rect -2500 1011 -2466 1013
rect -2242 1011 -2208 1013
rect -1800 1011 -1766 1013
rect -1542 1011 -1508 1013
rect -1100 1011 -1066 1013
rect -842 1011 -808 1013
rect -400 1011 -366 1013
rect -142 1011 -108 1013
rect 300 1011 334 1013
rect 558 1011 592 1013
rect 1000 1011 1034 1013
rect 1258 1011 1292 1013
rect 1700 1011 1734 1013
rect 1958 1011 1992 1013
rect 2400 1011 2434 1013
rect 2658 1011 2692 1013
rect 3100 1011 3134 1013
rect 3358 1011 3392 1013
rect 3800 1011 3834 1013
rect 4058 1011 4092 1013
rect -2500 981 -2466 983
rect -2242 981 -2208 983
rect -1800 981 -1766 983
rect -1542 981 -1508 983
rect -1100 981 -1066 983
rect -842 981 -808 983
rect -400 981 -366 983
rect -142 981 -108 983
rect 300 981 334 983
rect 558 981 592 983
rect 1000 981 1034 983
rect 1258 981 1292 983
rect 1700 981 1734 983
rect 1958 981 1992 983
rect 2400 981 2434 983
rect 2658 981 2692 983
rect 3100 981 3134 983
rect 3358 981 3392 983
rect 3800 981 3834 983
rect 4058 981 4092 983
rect -2500 947 -2466 949
rect -2242 947 -2208 949
rect -1800 947 -1766 949
rect -1542 947 -1508 949
rect -1100 947 -1066 949
rect -842 947 -808 949
rect -400 947 -366 949
rect -142 947 -108 949
rect 300 947 334 949
rect 558 947 592 949
rect 1000 947 1034 949
rect 1258 947 1292 949
rect 1700 947 1734 949
rect 1958 947 1992 949
rect 2400 947 2434 949
rect 2658 947 2692 949
rect 3100 947 3134 949
rect 3358 947 3392 949
rect 3800 947 3834 949
rect 4058 947 4092 949
rect -2500 943 -2466 945
rect -2242 943 -2208 945
rect -1800 943 -1766 945
rect -1542 943 -1508 945
rect -1100 943 -1066 945
rect -842 943 -808 945
rect -400 943 -366 945
rect -142 943 -108 945
rect 300 943 334 945
rect 558 943 592 945
rect 1000 943 1034 945
rect 1258 943 1292 945
rect 1700 943 1734 945
rect 1958 943 1992 945
rect 2400 943 2434 945
rect 2658 943 2692 945
rect 3100 943 3134 945
rect 3358 943 3392 945
rect 3800 943 3834 945
rect 4058 943 4092 945
rect -2500 909 -2466 911
rect -2242 909 -2208 911
rect -1800 909 -1766 911
rect -1542 909 -1508 911
rect -1100 909 -1066 911
rect -842 909 -808 911
rect -400 909 -366 911
rect -142 909 -108 911
rect 300 909 334 911
rect 558 909 592 911
rect 1000 909 1034 911
rect 1258 909 1292 911
rect 1700 909 1734 911
rect 1958 909 1992 911
rect 2400 909 2434 911
rect 2658 909 2692 911
rect 3100 909 3134 911
rect 3358 909 3392 911
rect 3800 909 3834 911
rect 4058 909 4092 911
rect -2500 875 -2466 877
rect -2242 875 -2208 877
rect -1800 875 -1766 877
rect -1542 875 -1508 877
rect -1100 875 -1066 877
rect -842 875 -808 877
rect -400 875 -366 877
rect -142 875 -108 877
rect 300 875 334 877
rect 558 875 592 877
rect 1000 875 1034 877
rect 1258 875 1292 877
rect 1700 875 1734 877
rect 1958 875 1992 877
rect 2400 875 2434 877
rect 2658 875 2692 877
rect 3100 875 3134 877
rect 3358 875 3392 877
rect 3800 875 3834 877
rect 4058 875 4092 877
rect -2500 837 -2466 839
rect -2242 837 -2208 839
rect -1800 837 -1766 839
rect -1542 837 -1508 839
rect -1100 837 -1066 839
rect -842 837 -808 839
rect -400 837 -366 839
rect -142 837 -108 839
rect 300 837 334 839
rect 558 837 592 839
rect 1000 837 1034 839
rect 1258 837 1292 839
rect 1700 837 1734 839
rect 1958 837 1992 839
rect 2400 837 2434 839
rect 2658 837 2692 839
rect 3100 837 3134 839
rect 3358 837 3392 839
rect 3800 837 3834 839
rect 4058 837 4092 839
rect -2500 807 -2466 809
rect -2242 807 -2208 809
rect -1800 807 -1766 809
rect -1542 807 -1508 809
rect -1100 807 -1066 809
rect -842 807 -808 809
rect -400 807 -366 809
rect -142 807 -108 809
rect 300 807 334 809
rect 558 807 592 809
rect 1000 807 1034 809
rect 1258 807 1292 809
rect 1700 807 1734 809
rect 1958 807 1992 809
rect 2400 807 2434 809
rect 2658 807 2692 809
rect 3100 807 3134 809
rect 3358 807 3392 809
rect 3800 807 3834 809
rect 4058 807 4092 809
rect -2500 803 -2466 805
rect -2242 803 -2208 805
rect -1800 803 -1766 805
rect -1542 803 -1508 805
rect -1100 803 -1066 805
rect -842 803 -808 805
rect -400 803 -366 805
rect -142 803 -108 805
rect 300 803 334 805
rect 558 803 592 805
rect 1000 803 1034 805
rect 1258 803 1292 805
rect 1700 803 1734 805
rect 1958 803 1992 805
rect 2400 803 2434 805
rect 2658 803 2692 805
rect 3100 803 3134 805
rect 3358 803 3392 805
rect 3800 803 3834 805
rect 4058 803 4092 805
rect -2500 765 -2466 767
rect -2242 765 -2208 767
rect -1800 765 -1766 767
rect -1542 765 -1508 767
rect -1100 765 -1066 767
rect -842 765 -808 767
rect -400 765 -366 767
rect -142 765 -108 767
rect 300 765 334 767
rect 558 765 592 767
rect 1000 765 1034 767
rect 1258 765 1292 767
rect 1700 765 1734 767
rect 1958 765 1992 767
rect 2400 765 2434 767
rect 2658 765 2692 767
rect 3100 765 3134 767
rect 3358 765 3392 767
rect 3800 765 3834 767
rect 4058 765 4092 767
rect -2500 739 -2466 741
rect -2242 739 -2208 741
rect -1800 739 -1766 741
rect -1542 739 -1508 741
rect -1100 739 -1066 741
rect -842 739 -808 741
rect -400 739 -366 741
rect -142 739 -108 741
rect 300 739 334 741
rect 558 739 592 741
rect 1000 739 1034 741
rect 1258 739 1292 741
rect 1700 739 1734 741
rect 1958 739 1992 741
rect 2400 739 2434 741
rect 2658 739 2692 741
rect 3100 739 3134 741
rect 3358 739 3392 741
rect 3800 739 3834 741
rect 4058 739 4092 741
rect -2500 731 -2466 733
rect -2242 731 -2208 733
rect -1800 731 -1766 733
rect -1542 731 -1508 733
rect -1100 731 -1066 733
rect -842 731 -808 733
rect -400 731 -366 733
rect -142 731 -108 733
rect 300 731 334 733
rect 558 731 592 733
rect 1000 731 1034 733
rect 1258 731 1292 733
rect 1700 731 1734 733
rect 1958 731 1992 733
rect 2400 731 2434 733
rect 2658 731 2692 733
rect 3100 731 3134 733
rect 3358 731 3392 733
rect 3800 731 3834 733
rect 4058 731 4092 733
rect -2500 693 -2466 695
rect -2242 693 -2208 695
rect -1800 693 -1766 695
rect -1542 693 -1508 695
rect -1100 693 -1066 695
rect -842 693 -808 695
rect -400 693 -366 695
rect -142 693 -108 695
rect 300 693 334 695
rect 558 693 592 695
rect 1000 693 1034 695
rect 1258 693 1292 695
rect 1700 693 1734 695
rect 1958 693 1992 695
rect 2400 693 2434 695
rect 2658 693 2692 695
rect 3100 693 3134 695
rect 3358 693 3392 695
rect 3800 693 3834 695
rect 4058 693 4092 695
rect -2500 671 -2466 673
rect -2242 671 -2208 673
rect -1800 671 -1766 673
rect -1542 671 -1508 673
rect -1100 671 -1066 673
rect -842 671 -808 673
rect -400 671 -366 673
rect -142 671 -108 673
rect 300 671 334 673
rect 558 671 592 673
rect 1000 671 1034 673
rect 1258 671 1292 673
rect 1700 671 1734 673
rect 1958 671 1992 673
rect 2400 671 2434 673
rect 2658 671 2692 673
rect 3100 671 3134 673
rect 3358 671 3392 673
rect 3800 671 3834 673
rect 4058 671 4092 673
rect -2500 659 -2466 661
rect -2242 659 -2208 661
rect -1800 659 -1766 661
rect -1542 659 -1508 661
rect -1100 659 -1066 661
rect -842 659 -808 661
rect -400 659 -366 661
rect -142 659 -108 661
rect 300 659 334 661
rect 558 659 592 661
rect 1000 659 1034 661
rect 1258 659 1292 661
rect 1700 659 1734 661
rect 1958 659 1992 661
rect 2400 659 2434 661
rect 2658 659 2692 661
rect 3100 659 3134 661
rect 3358 659 3392 661
rect 3800 659 3834 661
rect 4058 659 4092 661
rect -2500 621 -2466 623
rect -2242 621 -2208 623
rect -1800 621 -1766 623
rect -1542 621 -1508 623
rect -1100 621 -1066 623
rect -842 621 -808 623
rect -400 621 -366 623
rect -142 621 -108 623
rect 300 621 334 623
rect 558 621 592 623
rect 1000 621 1034 623
rect 1258 621 1292 623
rect 1700 621 1734 623
rect 1958 621 1992 623
rect 2400 621 2434 623
rect 2658 621 2692 623
rect 3100 621 3134 623
rect 3358 621 3392 623
rect 3800 621 3834 623
rect 4058 621 4092 623
rect -2500 603 -2466 605
rect -2242 603 -2208 605
rect -1800 603 -1766 605
rect -1542 603 -1508 605
rect -1100 603 -1066 605
rect -842 603 -808 605
rect -400 603 -366 605
rect -142 603 -108 605
rect 300 603 334 605
rect 558 603 592 605
rect 1000 603 1034 605
rect 1258 603 1292 605
rect 1700 603 1734 605
rect 1958 603 1992 605
rect 2400 603 2434 605
rect 2658 603 2692 605
rect 3100 603 3134 605
rect 3358 603 3392 605
rect 3800 603 3834 605
rect 4058 603 4092 605
rect -2500 587 -2466 589
rect -2242 587 -2208 589
rect -1800 587 -1766 589
rect -1542 587 -1508 589
rect -1100 587 -1066 589
rect -842 587 -808 589
rect -400 587 -366 589
rect -142 587 -108 589
rect 300 587 334 589
rect 558 587 592 589
rect 1000 587 1034 589
rect 1258 587 1292 589
rect 1700 587 1734 589
rect 1958 587 1992 589
rect 2400 587 2434 589
rect 2658 587 2692 589
rect 3100 587 3134 589
rect 3358 587 3392 589
rect 3800 587 3834 589
rect 4058 587 4092 589
rect -2500 549 -2466 551
rect -2242 549 -2208 551
rect -1800 549 -1766 551
rect -1542 549 -1508 551
rect -1100 549 -1066 551
rect -842 549 -808 551
rect -400 549 -366 551
rect -142 549 -108 551
rect 300 549 334 551
rect 558 549 592 551
rect 1000 549 1034 551
rect 1258 549 1292 551
rect 1700 549 1734 551
rect 1958 549 1992 551
rect 2400 549 2434 551
rect 2658 549 2692 551
rect 3100 549 3134 551
rect 3358 549 3392 551
rect 3800 549 3834 551
rect 4058 549 4092 551
rect -2500 535 -2466 537
rect -2242 535 -2208 537
rect -1800 535 -1766 537
rect -1542 535 -1508 537
rect -1100 535 -1066 537
rect -842 535 -808 537
rect -400 535 -366 537
rect -142 535 -108 537
rect 300 535 334 537
rect 558 535 592 537
rect 1000 535 1034 537
rect 1258 535 1292 537
rect 1700 535 1734 537
rect 1958 535 1992 537
rect 2400 535 2434 537
rect 2658 535 2692 537
rect 3100 535 3134 537
rect 3358 535 3392 537
rect 3800 535 3834 537
rect 4058 535 4092 537
rect -2500 515 -2466 517
rect -2242 515 -2208 517
rect -1800 515 -1766 517
rect -1542 515 -1508 517
rect -1100 515 -1066 517
rect -842 515 -808 517
rect -400 515 -366 517
rect -142 515 -108 517
rect 300 515 334 517
rect 558 515 592 517
rect 1000 515 1034 517
rect 1258 515 1292 517
rect 1700 515 1734 517
rect 1958 515 1992 517
rect 2400 515 2434 517
rect 2658 515 2692 517
rect 3100 515 3134 517
rect 3358 515 3392 517
rect 3800 515 3834 517
rect 4058 515 4092 517
rect -2500 477 -2466 479
rect -2242 477 -2208 479
rect -1800 477 -1766 479
rect -1542 477 -1508 479
rect -1100 477 -1066 479
rect -842 477 -808 479
rect -400 477 -366 479
rect -142 477 -108 479
rect 300 477 334 479
rect 558 477 592 479
rect 1000 477 1034 479
rect 1258 477 1292 479
rect 1700 477 1734 479
rect 1958 477 1992 479
rect 2400 477 2434 479
rect 2658 477 2692 479
rect 3100 477 3134 479
rect 3358 477 3392 479
rect 3800 477 3834 479
rect 4058 477 4092 479
rect -2500 467 -2466 469
rect -2242 467 -2208 469
rect -1800 467 -1766 469
rect -1542 467 -1508 469
rect -1100 467 -1066 469
rect -842 467 -808 469
rect -400 467 -366 469
rect -142 467 -108 469
rect 300 467 334 469
rect 558 467 592 469
rect 1000 467 1034 469
rect 1258 467 1292 469
rect 1700 467 1734 469
rect 1958 467 1992 469
rect 2400 467 2434 469
rect 2658 467 2692 469
rect 3100 467 3134 469
rect 3358 467 3392 469
rect 3800 467 3834 469
rect 4058 467 4092 469
rect -2500 443 -2466 445
rect -2242 443 -2208 445
rect -1800 443 -1766 445
rect -1542 443 -1508 445
rect -1100 443 -1066 445
rect -842 443 -808 445
rect -400 443 -366 445
rect -142 443 -108 445
rect 300 443 334 445
rect 558 443 592 445
rect 1000 443 1034 445
rect 1258 443 1292 445
rect 1700 443 1734 445
rect 1958 443 1992 445
rect 2400 443 2434 445
rect 2658 443 2692 445
rect 3100 443 3134 445
rect 3358 443 3392 445
rect 3800 443 3834 445
rect 4058 443 4092 445
rect -2500 405 -2466 407
rect -2242 405 -2208 407
rect -1800 405 -1766 407
rect -1542 405 -1508 407
rect -1100 405 -1066 407
rect -842 405 -808 407
rect -400 405 -366 407
rect -142 405 -108 407
rect 300 405 334 407
rect 558 405 592 407
rect 1000 405 1034 407
rect 1258 405 1292 407
rect 1700 405 1734 407
rect 1958 405 1992 407
rect 2400 405 2434 407
rect 2658 405 2692 407
rect 3100 405 3134 407
rect 3358 405 3392 407
rect 3800 405 3834 407
rect 4058 405 4092 407
rect -2500 399 -2466 401
rect -2242 399 -2208 401
rect -1800 399 -1766 401
rect -1542 399 -1508 401
rect -1100 399 -1066 401
rect -842 399 -808 401
rect -400 399 -366 401
rect -142 399 -108 401
rect 300 399 334 401
rect 558 399 592 401
rect 1000 399 1034 401
rect 1258 399 1292 401
rect 1700 399 1734 401
rect 1958 399 1992 401
rect 2400 399 2434 401
rect 2658 399 2692 401
rect 3100 399 3134 401
rect 3358 399 3392 401
rect 3800 399 3834 401
rect 4058 399 4092 401
rect -2500 371 -2466 373
rect -2242 371 -2208 373
rect -1800 371 -1766 373
rect -1542 371 -1508 373
rect -1100 371 -1066 373
rect -842 371 -808 373
rect -400 371 -366 373
rect -142 371 -108 373
rect 300 371 334 373
rect 558 371 592 373
rect 1000 371 1034 373
rect 1258 371 1292 373
rect 1700 371 1734 373
rect 1958 371 1992 373
rect 2400 371 2434 373
rect 2658 371 2692 373
rect 3100 371 3134 373
rect 3358 371 3392 373
rect 3800 371 3834 373
rect 4058 371 4092 373
rect -2500 331 -2466 335
rect -2242 331 -2208 335
rect -1800 331 -1766 335
rect -1542 331 -1508 335
rect -1100 331 -1066 335
rect -842 331 -808 335
rect -400 331 -366 335
rect -142 331 -108 335
rect 300 331 334 335
rect 558 331 592 335
rect 1000 331 1034 335
rect 1258 331 1292 335
rect 1700 331 1734 335
rect 1958 331 1992 335
rect 2400 331 2434 335
rect 2658 331 2692 335
rect 3100 331 3134 335
rect 3358 331 3392 335
rect 3800 331 3834 335
rect 4058 331 4092 335
rect -2500 299 -2466 301
rect -2242 299 -2208 301
rect -1800 299 -1766 301
rect -1542 299 -1508 301
rect -1100 299 -1066 301
rect -842 299 -808 301
rect -400 299 -366 301
rect -142 299 -108 301
rect 300 299 334 301
rect 558 299 592 301
rect 1000 299 1034 301
rect 1258 299 1292 301
rect 1700 299 1734 301
rect 1958 299 1992 301
rect 2400 299 2434 301
rect 2658 299 2692 301
rect 3100 299 3134 301
rect 3358 299 3392 301
rect 3800 299 3834 301
rect 4058 299 4092 301
rect -2500 261 -2466 265
rect -2242 261 -2208 265
rect -1800 261 -1766 265
rect -1542 261 -1508 265
rect -1100 261 -1066 265
rect -842 261 -808 265
rect -400 261 -366 265
rect -142 261 -108 265
rect 300 261 334 265
rect 558 261 592 265
rect 1000 261 1034 265
rect 1258 261 1292 265
rect 1700 261 1734 265
rect 1958 261 1992 265
rect 2400 261 2434 265
rect 2658 261 2692 265
rect 3100 261 3134 265
rect 3358 261 3392 265
rect 3800 261 3834 265
rect 4058 261 4092 265
rect -2500 227 -2466 229
rect -2242 227 -2208 229
rect -1800 227 -1766 229
rect -1542 227 -1508 229
rect -1100 227 -1066 229
rect -842 227 -808 229
rect -400 227 -366 229
rect -142 227 -108 229
rect 300 227 334 229
rect 558 227 592 229
rect 1000 227 1034 229
rect 1258 227 1292 229
rect 1700 227 1734 229
rect 1958 227 1992 229
rect 2400 227 2434 229
rect 2658 227 2692 229
rect 3100 227 3134 229
rect 3358 227 3392 229
rect 3800 227 3834 229
rect 4058 227 4092 229
rect -2500 195 -2466 197
rect -2242 195 -2208 197
rect -1800 195 -1766 197
rect -1542 195 -1508 197
rect -1100 195 -1066 197
rect -842 195 -808 197
rect -400 195 -366 197
rect -142 195 -108 197
rect 300 195 334 197
rect 558 195 592 197
rect 1000 195 1034 197
rect 1258 195 1292 197
rect 1700 195 1734 197
rect 1958 195 1992 197
rect 2400 195 2434 197
rect 2658 195 2692 197
rect 3100 195 3134 197
rect 3358 195 3392 197
rect 3800 195 3834 197
rect 4058 195 4092 197
rect -2500 189 -2466 191
rect -2242 189 -2208 191
rect -1800 189 -1766 191
rect -1542 189 -1508 191
rect -1100 189 -1066 191
rect -842 189 -808 191
rect -400 189 -366 191
rect -142 189 -108 191
rect 300 189 334 191
rect 558 189 592 191
rect 1000 189 1034 191
rect 1258 189 1292 191
rect 1700 189 1734 191
rect 1958 189 1992 191
rect 2400 189 2434 191
rect 2658 189 2692 191
rect 3100 189 3134 191
rect 3358 189 3392 191
rect 3800 189 3834 191
rect 4058 189 4092 191
rect -2500 155 -2466 157
rect -2242 155 -2208 157
rect -1800 155 -1766 157
rect -1542 155 -1508 157
rect -1100 155 -1066 157
rect -842 155 -808 157
rect -400 155 -366 157
rect -142 155 -108 157
rect 300 155 334 157
rect 558 155 592 157
rect 1000 155 1034 157
rect 1258 155 1292 157
rect 1700 155 1734 157
rect 1958 155 1992 157
rect 2400 155 2434 157
rect 2658 155 2692 157
rect 3100 155 3134 157
rect 3358 155 3392 157
rect 3800 155 3834 157
rect 4058 155 4092 157
rect -2500 127 -2466 129
rect -2242 127 -2208 129
rect -1800 127 -1766 129
rect -1542 127 -1508 129
rect -1100 127 -1066 129
rect -842 127 -808 129
rect -400 127 -366 129
rect -142 127 -108 129
rect 300 127 334 129
rect 558 127 592 129
rect 1000 127 1034 129
rect 1258 127 1292 129
rect 1700 127 1734 129
rect 1958 127 1992 129
rect 2400 127 2434 129
rect 2658 127 2692 129
rect 3100 127 3134 129
rect 3358 127 3392 129
rect 3800 127 3834 129
rect 4058 127 4092 129
rect -2500 117 -2466 119
rect -2242 117 -2208 119
rect -1800 117 -1766 119
rect -1542 117 -1508 119
rect -1100 117 -1066 119
rect -842 117 -808 119
rect -400 117 -366 119
rect -142 117 -108 119
rect 300 117 334 119
rect 558 117 592 119
rect 1000 117 1034 119
rect 1258 117 1292 119
rect 1700 117 1734 119
rect 1958 117 1992 119
rect 2400 117 2434 119
rect 2658 117 2692 119
rect 3100 117 3134 119
rect 3358 117 3392 119
rect 3800 117 3834 119
rect 4058 117 4092 119
rect -2500 83 -2466 85
rect -2242 83 -2208 85
rect -1800 83 -1766 85
rect -1542 83 -1508 85
rect -1100 83 -1066 85
rect -842 83 -808 85
rect -400 83 -366 85
rect -142 83 -108 85
rect 300 83 334 85
rect 558 83 592 85
rect 1000 83 1034 85
rect 1258 83 1292 85
rect 1700 83 1734 85
rect 1958 83 1992 85
rect 2400 83 2434 85
rect 2658 83 2692 85
rect 3100 83 3134 85
rect 3358 83 3392 85
rect 3800 83 3834 85
rect 4058 83 4092 85
rect -2500 59 -2466 61
rect -2242 59 -2208 61
rect -1800 59 -1766 61
rect -1542 59 -1508 61
rect -1100 59 -1066 61
rect -842 59 -808 61
rect -400 59 -366 61
rect -142 59 -108 61
rect 300 59 334 61
rect 558 59 592 61
rect 1000 59 1034 61
rect 1258 59 1292 61
rect 1700 59 1734 61
rect 1958 59 1992 61
rect 2400 59 2434 61
rect 2658 59 2692 61
rect 3100 59 3134 61
rect 3358 59 3392 61
rect 3800 59 3834 61
rect 4058 59 4092 61
rect -2500 45 -2466 47
rect -2242 45 -2208 47
rect -1800 45 -1766 47
rect -1542 45 -1508 47
rect -1100 45 -1066 47
rect -842 45 -808 47
rect -400 45 -366 47
rect -142 45 -108 47
rect 300 45 334 47
rect 558 45 592 47
rect 1000 45 1034 47
rect 1258 45 1292 47
rect 1700 45 1734 47
rect 1958 45 1992 47
rect 2400 45 2434 47
rect 2658 45 2692 47
rect 3100 45 3134 47
rect 3358 45 3392 47
rect 3800 45 3834 47
rect 4058 45 4092 47
rect -2500 11 -2466 13
rect -2242 11 -2208 13
rect -1800 11 -1766 13
rect -1542 11 -1508 13
rect -1100 11 -1066 13
rect -842 11 -808 13
rect -400 11 -366 13
rect -142 11 -108 13
rect 300 11 334 13
rect 558 11 592 13
rect 1000 11 1034 13
rect 1258 11 1292 13
rect 1700 11 1734 13
rect 1958 11 1992 13
rect 2400 11 2434 13
rect 2658 11 2692 13
rect 3100 11 3134 13
rect 3358 11 3392 13
rect 3800 11 3834 13
rect 4058 11 4092 13
rect -2500 -9 -2466 -7
rect -2242 -9 -2208 -7
rect -1800 -9 -1766 -7
rect -1542 -9 -1508 -7
rect -1100 -9 -1066 -7
rect -842 -9 -808 -7
rect -400 -9 -366 -7
rect -142 -9 -108 -7
rect 300 -9 334 -7
rect 558 -9 592 -7
rect 1000 -9 1034 -7
rect 1258 -9 1292 -7
rect 1700 -9 1734 -7
rect 1958 -9 1992 -7
rect 2400 -9 2434 -7
rect 2658 -9 2692 -7
rect 3100 -9 3134 -7
rect 3358 -9 3392 -7
rect 3800 -9 3834 -7
rect 4058 -9 4092 -7
rect -2500 -27 -2466 -25
rect -2242 -27 -2208 -25
rect -1800 -27 -1766 -25
rect -1542 -27 -1508 -25
rect -1100 -27 -1066 -25
rect -842 -27 -808 -25
rect -400 -27 -366 -25
rect -142 -27 -108 -25
rect 300 -27 334 -25
rect 558 -27 592 -25
rect 1000 -27 1034 -25
rect 1258 -27 1292 -25
rect 1700 -27 1734 -25
rect 1958 -27 1992 -25
rect 2400 -27 2434 -25
rect 2658 -27 2692 -25
rect 3100 -27 3134 -25
rect 3358 -27 3392 -25
rect 3800 -27 3834 -25
rect 4058 -27 4092 -25
rect -2374 -179 -2372 -145
rect -2338 -179 -2334 -145
rect -1674 -179 -1672 -145
rect -1638 -179 -1634 -145
rect -974 -179 -972 -145
rect -938 -179 -934 -145
rect -274 -179 -272 -145
rect -238 -179 -234 -145
rect 426 -179 428 -145
rect 462 -179 466 -145
rect 1126 -179 1128 -145
rect 1162 -179 1166 -145
rect 1826 -179 1828 -145
rect 1862 -179 1866 -145
rect 2526 -179 2528 -145
rect 2562 -179 2566 -145
rect 3226 -179 3228 -145
rect 3262 -179 3266 -145
rect 3926 -179 3928 -145
rect 3962 -179 3966 -145
<< metal1 >>
rect -2642 2443 3794 2603
rect -2202 -817 4234 -657
<< metal2 >>
rect -2712 2116 4043 2216
rect -2427 -323 4027 -238
use nfet_w10_l1  nfet_w10_l1_0
array 0 9 700 0 0 0
timestamp 1635946216
transform 1 0 372 0 1 99
box -3014 -756 -2438 2344
<< end >>
