magic
tech sky130A
magscale 1 4
timestamp 1632393576
<< pwell >>
rect -619 -1874 619 1874
<< nmos >>
rect -226 1054 -154 1454
rect -36 1054 36 1454
rect 154 1054 226 1454
rect -226 218 -154 618
rect -36 218 36 618
rect 154 218 226 618
rect -226 -618 -154 -218
rect -36 -618 36 -218
rect 154 -618 226 -218
rect -226 -1454 -154 -1054
rect -36 -1454 36 -1054
rect 154 -1454 226 -1054
<< ndiff >>
rect -343 1430 -226 1454
rect -343 1078 -319 1430
rect -251 1078 -226 1430
rect -343 1054 -226 1078
rect -154 1430 -36 1454
rect -154 1078 -129 1430
rect -61 1078 -36 1430
rect -154 1054 -36 1078
rect 36 1430 154 1454
rect 36 1078 61 1430
rect 129 1078 154 1430
rect 36 1054 154 1078
rect 226 1430 343 1454
rect 226 1078 251 1430
rect 319 1078 343 1430
rect 226 1054 343 1078
rect -343 594 -226 618
rect -343 242 -319 594
rect -251 242 -226 594
rect -343 218 -226 242
rect -154 594 -36 618
rect -154 242 -129 594
rect -61 242 -36 594
rect -154 218 -36 242
rect 36 594 154 618
rect 36 242 61 594
rect 129 242 154 594
rect 36 218 154 242
rect 226 594 343 618
rect 226 242 251 594
rect 319 242 343 594
rect 226 218 343 242
rect -343 -242 -226 -218
rect -343 -594 -319 -242
rect -251 -594 -226 -242
rect -343 -618 -226 -594
rect -154 -242 -36 -218
rect -154 -594 -129 -242
rect -61 -594 -36 -242
rect -154 -618 -36 -594
rect 36 -242 154 -218
rect 36 -594 61 -242
rect 129 -594 154 -242
rect 36 -618 154 -594
rect 226 -242 343 -218
rect 226 -594 251 -242
rect 319 -594 343 -242
rect 226 -618 343 -594
rect -343 -1078 -226 -1054
rect -343 -1430 -319 -1078
rect -251 -1430 -226 -1078
rect -343 -1454 -226 -1430
rect -154 -1078 -36 -1054
rect -154 -1430 -129 -1078
rect -61 -1430 -36 -1078
rect -154 -1454 -36 -1430
rect 36 -1078 154 -1054
rect 36 -1430 61 -1078
rect 129 -1430 154 -1078
rect 36 -1454 154 -1430
rect 226 -1078 343 -1054
rect 226 -1430 251 -1078
rect 319 -1430 343 -1078
rect 226 -1454 343 -1430
<< ndiffc >>
rect -319 1078 -251 1430
rect -129 1078 -61 1430
rect 61 1078 129 1430
rect 251 1078 319 1430
rect -319 242 -251 594
rect -129 242 -61 594
rect 61 242 129 594
rect 251 242 319 594
rect -319 -594 -251 -242
rect -129 -594 -61 -242
rect 61 -594 129 -242
rect 251 -594 319 -242
rect -319 -1430 -251 -1078
rect -129 -1430 -61 -1078
rect 61 -1430 129 -1078
rect 251 -1430 319 -1078
<< psubdiff >>
rect -547 1734 -355 1802
rect 355 1734 547 1802
rect -547 1610 -479 1734
rect 479 1610 547 1734
rect -547 -1734 -479 -1610
rect 479 -1734 547 -1610
rect -547 -1802 -355 -1734
rect 355 -1802 547 -1734
<< psubdiffcont >>
rect -355 1734 355 1802
rect -547 -1610 -479 1610
rect 479 -1610 547 1610
rect -355 -1802 355 -1734
<< poly >>
rect -256 1598 -124 1630
rect -256 1530 -224 1598
rect -156 1530 -124 1598
rect -256 1498 -124 1530
rect 124 1598 256 1630
rect 124 1530 156 1598
rect 224 1530 256 1598
rect -226 1454 -154 1498
rect -36 1454 36 1506
rect 124 1498 256 1530
rect 154 1454 226 1498
rect -226 1002 -154 1054
rect -36 1010 36 1054
rect -66 978 66 1010
rect 154 1002 226 1054
rect -66 910 -34 978
rect 34 910 66 978
rect -66 878 66 910
rect -66 762 66 794
rect -66 694 -34 762
rect 34 694 66 762
rect -226 618 -154 670
rect -66 662 66 694
rect -36 618 36 662
rect 154 618 226 670
rect -226 174 -154 218
rect -256 142 -124 174
rect -36 166 36 218
rect 154 174 226 218
rect -256 74 -224 142
rect -156 74 -124 142
rect -256 42 -124 74
rect 124 142 256 174
rect 124 74 156 142
rect 224 74 256 142
rect 124 42 256 74
rect -256 -74 -124 -42
rect -256 -142 -224 -74
rect -156 -142 -124 -74
rect -256 -174 -124 -142
rect 124 -74 256 -42
rect 124 -142 156 -74
rect 224 -142 256 -74
rect -226 -218 -154 -174
rect -36 -218 36 -166
rect 124 -174 256 -142
rect 154 -218 226 -174
rect -226 -670 -154 -618
rect -36 -662 36 -618
rect -66 -694 66 -662
rect 154 -670 226 -618
rect -66 -762 -34 -694
rect 34 -762 66 -694
rect -66 -794 66 -762
rect -66 -910 66 -878
rect -66 -978 -34 -910
rect 34 -978 66 -910
rect -226 -1054 -154 -1002
rect -66 -1010 66 -978
rect -36 -1054 36 -1010
rect 154 -1054 226 -1002
rect -226 -1498 -154 -1454
rect -256 -1530 -124 -1498
rect -36 -1506 36 -1454
rect 154 -1498 226 -1454
rect -256 -1598 -224 -1530
rect -156 -1598 -124 -1530
rect -256 -1630 -124 -1598
rect 124 -1530 256 -1498
rect 124 -1598 156 -1530
rect 224 -1598 256 -1530
rect 124 -1630 256 -1598
<< polycont >>
rect -224 1530 -156 1598
rect 156 1530 224 1598
rect -34 910 34 978
rect -34 694 34 762
rect -224 74 -156 142
rect 156 74 224 142
rect -224 -142 -156 -74
rect 156 -142 224 -74
rect -34 -762 34 -694
rect -34 -978 34 -910
rect -224 -1598 -156 -1530
rect 156 -1598 224 -1530
<< locali >>
rect -547 1734 -355 1802
rect 355 1734 547 1802
rect -547 1610 -479 1734
rect 479 1610 547 1734
rect -256 1530 -224 1598
rect -156 1530 -124 1598
rect 124 1530 156 1598
rect 224 1530 256 1598
rect -319 1430 -251 1462
rect -319 1046 -251 1078
rect -129 1430 -61 1462
rect -129 1046 -61 1078
rect 61 1430 129 1462
rect 61 1046 129 1078
rect 251 1430 319 1462
rect 251 1046 319 1078
rect -66 910 -34 978
rect 34 910 66 978
rect -66 694 -34 762
rect 34 694 66 762
rect -319 594 -251 626
rect -319 210 -251 242
rect -129 594 -61 626
rect -129 210 -61 242
rect 61 594 129 626
rect 61 210 129 242
rect 251 594 319 626
rect 251 210 319 242
rect -256 74 -224 142
rect -156 74 -124 142
rect 124 74 156 142
rect 224 74 256 142
rect -256 -142 -224 -74
rect -156 -142 -124 -74
rect 124 -142 156 -74
rect 224 -142 256 -74
rect -319 -242 -251 -210
rect -319 -626 -251 -594
rect -129 -242 -61 -210
rect -129 -626 -61 -594
rect 61 -242 129 -210
rect 61 -626 129 -594
rect 251 -242 319 -210
rect 251 -626 319 -594
rect -66 -762 -34 -694
rect 34 -762 66 -694
rect -66 -978 -34 -910
rect 34 -978 66 -910
rect -319 -1078 -251 -1046
rect -319 -1462 -251 -1430
rect -129 -1078 -61 -1046
rect -129 -1462 -61 -1430
rect 61 -1078 129 -1046
rect 61 -1462 129 -1430
rect 251 -1078 319 -1046
rect 251 -1462 319 -1430
rect -256 -1598 -224 -1530
rect -156 -1598 -124 -1530
rect 124 -1598 156 -1530
rect 224 -1598 256 -1530
rect -547 -1734 -479 -1610
rect 479 -1734 547 -1610
rect -547 -1802 -355 -1734
rect 355 -1802 547 -1734
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -513 -1768 513 1768
string parameters w 1 l 0.18 m 4 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
