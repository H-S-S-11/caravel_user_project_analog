* SPICE3 file created from diffamp.ext - technology: sky130A

X0 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 VOPAMP VOP ISINK VGND sky130_fd_pr__nfet_01v8 ad=-0p pd=0u as=-0p ps=0u w=1e+06u l=180000u
X2 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X3 VONAMP VON ISINK VGND sky130_fd_pr__nfet_01v8 ad=-0p pd=0u as=-0p ps=0u w=1e+06u l=180000u
X4 VGND VONAMP ISINK VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=-0p ps=0u w=1e+06u l=180000u
X5 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X6 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X7 VONAMP VONAMP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=-0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X8 VPWR VONAMP VOPAMP VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=1e+06u l=180000u
X9 VPWR VONAMP VONAMP VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=1e+06u l=180000u
X10 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X11 VOPAMP VONAMP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=-0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X12 VPWR VONAMP VONAMP VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=1e+06u l=180000u
X13 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X14 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X15 VPWR VONAMP VOPAMP VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=1e+06u l=180000u
X16 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X17 VPWR VOPAMP VOUT VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 VGND VOPAMP VOUT VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 VPWR VGND 11.52fF
C1 VONAMP VGND 2.51fF
