magic
tech sky130A
timestamp 1633982189
<< nsonos >>
rect -7 -50 9 50
<< ndiff >>
rect -52 40 -7 50
rect -52 -40 -42 40
rect -22 -40 -7 40
rect -52 -50 -7 -40
rect 9 40 58 50
rect 9 -40 28 40
rect 48 -40 58 40
rect 9 -50 58 -40
<< ndiffc >>
rect -42 -40 -22 40
rect 28 -40 48 40
<< psubdiff >>
rect -102 130 108 150
rect -102 -120 -82 130
rect 88 -120 108 130
rect -102 -140 -42 -120
rect 48 -140 108 -120
<< psubdiffcont >>
rect -42 -140 48 -120
<< poly >>
rect -22 100 28 110
rect -22 80 -12 100
rect 18 80 28 100
rect -22 70 28 80
rect -7 50 9 70
rect -7 -70 9 -50
<< polycont >>
rect -12 80 18 100
<< locali >>
rect -22 100 28 110
rect -22 80 -12 100
rect 18 80 28 100
rect -22 70 28 80
rect -52 40 -22 50
rect -52 -40 -42 40
rect -52 -50 -22 -40
rect 28 40 58 50
rect 48 -40 58 40
rect 28 -50 58 -40
rect -52 -140 -42 -120
rect 48 -140 58 -120
<< properties >>
string gencell sky130_fd_bs_flash__special_sonosfet_star
string FIXED_BBOX -82 -130 82 130
string parameters w 1 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
