magic
tech sky130A
magscale 1 2
timestamp 1632652117
<< locali >>
rect 1760 1900 1860 1920
rect 1760 1840 1780 1900
rect 1840 1840 1860 1900
rect 1760 1540 1860 1840
rect 1760 1480 1780 1540
rect 1840 1480 1860 1540
rect 1760 1460 1860 1480
<< viali >>
rect 1780 1840 1840 1900
rect 1780 1480 1840 1540
<< metal1 >>
rect -240 2420 40 2800
rect 480 2180 1620 2800
rect 2060 2460 2400 2800
rect 2720 2680 4420 2800
rect 2720 2600 3620 2680
rect 1140 1980 1620 2180
rect 4040 2120 4420 2680
rect 4560 2080 4660 2800
rect 4940 2140 5360 2800
rect -440 1900 1860 1920
rect -440 1840 1780 1900
rect 1840 1840 1860 1900
rect -440 1820 1860 1840
rect 2900 1780 3900 1880
rect 460 1640 2000 1740
rect 460 1420 580 1640
rect 1760 1540 1860 1560
rect 1760 1480 1780 1540
rect 1840 1480 1860 1540
rect 1230 1380 1600 1470
rect -440 1270 540 1350
rect 1500 1340 1600 1380
rect 1760 1340 1860 1480
rect 1500 1240 1860 1340
rect 1900 1320 2000 1640
rect 3800 1280 3900 1780
rect -440 1160 540 1240
rect 460 860 580 1080
rect 1900 860 2000 1220
rect 460 760 2000 860
rect 3800 720 3900 840
rect 2880 620 3900 720
use preamp  preamp_0
timestamp 1632332974
transform 1 0 -145 0 1 115
box -255 -115 1909 2460
use decision  decision_0
timestamp 1632485541
transform 1 0 2020 0 1 145
box -120 -245 1711 2620
use diffamp  diffamp_0
timestamp 1632488633
transform 1 0 4840 0 1 -1080
box -940 980 620 3400
<< labels >>
rlabel metal1 -440 1270 -430 1350 1 VP
port 2 n
rlabel metal1 -440 1160 -430 1240 1 VN
port 1 n
rlabel metal1 480 2760 1620 2800 1 VGND
port 5 n
rlabel metal1 2720 2760 4420 2800 1 VGND
port 5 n
rlabel metal1 -440 1820 -420 1920 1 BIASN
port 3 n
rlabel metal1 4560 2760 4660 2800 1 VOUT
port 6 n
rlabel metal1 4940 2760 5360 2800 1 VDD1v8
port 7 n
rlabel metal1 2060 2760 2400 2800 1 VDD3v3
port 4 n
rlabel metal1 -240 2760 40 2800 1 VDD3v3
port 4 n
<< end >>
